VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 221.8 BY 370.6 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  185.8 54.4 186.6 55.2 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  207.6 54.4 208.4 55.2 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  70.2 299.2 71.0 300.0 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  70.2 321.2 71.0 322.0 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  70.2 339.2 71.0 340.0 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  70.2 361.2 71.0 362.0 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  7.6 8.6 8.4 9.4 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  7.6 30.6 8.4 31.4 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  51.1 0.0 51.7 9.8 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  192.4 117.6 193.2 120.6 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  199.2 117.6 200.0 120.6 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  144.7 348.0 145.5 348.8 ;
         LAYER m3 ;
         RECT  201.7 243.7 202.3 244.3 ;
         LAYER m3 ;
         RECT  210.5 65.4 211.3 66.2 ;
         LAYER m3 ;
         RECT  208.5 285.3 209.1 285.9 ;
         LAYER m3 ;
         RECT  208.5 326.9 209.1 327.5 ;
         LAYER m3 ;
         RECT  118.7 223.2 119.5 224.0 ;
         LAYER m3 ;
         RECT  188.0 264.4 188.8 265.2 ;
         LAYER m3 ;
         RECT  194.9 222.9 195.5 223.5 ;
         LAYER m3 ;
         RECT  188.0 181.2 188.8 182.0 ;
         LAYER m3 ;
         RECT  181.3 181.3 181.9 181.9 ;
         LAYER m3 ;
         RECT  103.7 202.4 104.5 203.2 ;
         LAYER m3 ;
         RECT  208.5 264.5 209.1 265.1 ;
         LAYER m3 ;
         RECT  201.7 326.9 202.3 327.5 ;
         LAYER m3 ;
         RECT  194.9 326.9 195.5 327.5 ;
         LAYER m3 ;
         RECT  188.0 368.4 188.8 369.2 ;
         LAYER m3 ;
         RECT  165.5 244.0 166.3 244.8 ;
         LAYER m3 ;
         RECT  194.9 285.3 195.5 285.9 ;
         LAYER m3 ;
         RECT  194.6 160.8 195.4 161.6 ;
         LAYER m3 ;
         RECT  12.4 263.2 13.2 264.0 ;
         LAYER m3 ;
         RECT  103.7 223.2 104.5 224.0 ;
         LAYER m3 ;
         RECT  208.5 306.1 209.1 306.7 ;
         LAYER m3 ;
         RECT  194.9 347.7 195.5 348.3 ;
         LAYER m3 ;
         RECT  188.0 285.2 188.8 286.0 ;
         LAYER m3 ;
         RECT  195.6 79.0 196.4 79.8 ;
         LAYER m3 ;
         RECT  12.4 196.0 13.2 196.8 ;
         LAYER m3 ;
         RECT  181.3 285.3 181.9 285.9 ;
         LAYER m3 ;
         RECT  18.8 240.8 19.6 241.6 ;
         LAYER m3 ;
         RECT  201.7 306.1 202.3 306.7 ;
         LAYER m3 ;
         RECT  6.0 263.2 6.8 264.0 ;
         LAYER m3 ;
         RECT  201.7 264.5 202.3 265.1 ;
         LAYER m3 ;
         RECT  144.7 223.2 145.5 224.0 ;
         LAYER m3 ;
         RECT  12.4 218.4 13.2 219.2 ;
         LAYER m3 ;
         RECT  208.5 181.3 209.1 181.9 ;
         LAYER m3 ;
         RECT  144.7 244.0 145.5 244.8 ;
         LAYER m3 ;
         RECT  6.0 196.0 6.8 196.8 ;
         LAYER m3 ;
         RECT  82.6 99.6 83.4 100.4 ;
         LAYER m3 ;
         RECT  165.5 348.0 166.3 348.8 ;
         LAYER m3 ;
         RECT  144.7 327.2 145.5 328.0 ;
         LAYER m3 ;
         RECT  201.4 160.8 202.2 161.6 ;
         LAYER m3 ;
         RECT  -0.4 19.6 0.4 20.4 ;
         LAYER m3 ;
         RECT  165.5 306.4 166.3 307.2 ;
         LAYER m3 ;
         RECT  165.5 327.2 166.3 328.0 ;
         LAYER m3 ;
         RECT  187.8 160.8 188.6 161.6 ;
         LAYER m3 ;
         RECT  165.5 285.6 166.3 286.4 ;
         LAYER m3 ;
         RECT  188.7 65.4 189.5 66.2 ;
         LAYER m3 ;
         RECT  165.5 202.4 166.3 203.2 ;
         LAYER m3 ;
         RECT  12.4 240.8 13.2 241.6 ;
         LAYER m3 ;
         RECT  73.1 350.2 73.9 351.0 ;
         LAYER m3 ;
         RECT  204.0 130.4 204.8 131.2 ;
         LAYER m3 ;
         RECT  6.0 240.8 6.8 241.6 ;
         LAYER m3 ;
         RECT  201.7 181.3 202.3 181.9 ;
         LAYER m3 ;
         RECT  103.7 264.8 104.5 265.6 ;
         LAYER m3 ;
         RECT  202.4 79.0 203.2 79.8 ;
         LAYER m3 ;
         RECT  194.9 264.5 195.5 265.1 ;
         LAYER m3 ;
         RECT  144.7 264.8 145.5 265.6 ;
         LAYER m3 ;
         RECT  194.9 368.5 195.5 369.1 ;
         LAYER m3 ;
         RECT  118.7 264.8 119.5 265.6 ;
         LAYER m3 ;
         RECT  194.9 306.1 195.5 306.7 ;
         LAYER m3 ;
         RECT  181.3 202.1 181.9 202.7 ;
         LAYER m3 ;
         RECT  181.3 222.9 181.9 223.5 ;
         LAYER m3 ;
         RECT  188.0 222.8 188.8 223.6 ;
         LAYER m3 ;
         RECT  194.9 181.3 195.5 181.9 ;
         LAYER m3 ;
         RECT  73.1 310.2 73.9 311.0 ;
         LAYER m3 ;
         RECT  194.9 243.7 195.5 244.3 ;
         LAYER m3 ;
         RECT  188.0 347.6 188.8 348.4 ;
         LAYER m3 ;
         RECT  208.5 347.7 209.1 348.3 ;
         LAYER m3 ;
         RECT  6.0 173.6 6.8 174.4 ;
         LAYER m3 ;
         RECT  165.5 264.8 166.3 265.6 ;
         LAYER m3 ;
         RECT  82.6 59.6 83.4 60.4 ;
         LAYER m3 ;
         RECT  165.5 223.2 166.3 224.0 ;
         LAYER m3 ;
         RECT  201.7 222.9 202.3 223.5 ;
         LAYER m3 ;
         RECT  82.6 139.6 83.4 140.4 ;
         LAYER m3 ;
         RECT  201.7 202.1 202.3 202.7 ;
         LAYER m3 ;
         RECT  181.3 264.5 181.9 265.1 ;
         LAYER m3 ;
         RECT  18.8 263.2 19.6 264.0 ;
         LAYER m3 ;
         RECT  18.8 173.6 19.6 174.4 ;
         LAYER m3 ;
         RECT  201.7 347.7 202.3 348.3 ;
         LAYER m3 ;
         RECT  195.0 96.4 195.8 97.2 ;
         LAYER m3 ;
         RECT  201.8 96.4 202.6 97.2 ;
         LAYER m3 ;
         RECT  201.7 368.5 202.3 369.1 ;
         LAYER m3 ;
         RECT  188.0 202.0 188.8 202.8 ;
         LAYER m3 ;
         RECT  18.8 196.0 19.6 196.8 ;
         LAYER m3 ;
         RECT  82.6 19.6 83.4 20.4 ;
         LAYER m3 ;
         RECT  194.9 202.1 195.5 202.7 ;
         LAYER m3 ;
         RECT  188.0 306.0 188.8 306.8 ;
         LAYER m3 ;
         RECT  103.7 244.0 104.5 244.8 ;
         LAYER m3 ;
         RECT  118.7 244.0 119.5 244.8 ;
         LAYER m3 ;
         RECT  144.7 202.4 145.5 203.2 ;
         LAYER m3 ;
         RECT  144.7 306.4 145.5 307.2 ;
         LAYER m3 ;
         RECT  197.2 130.4 198.0 131.2 ;
         LAYER m3 ;
         RECT  208.5 368.5 209.1 369.1 ;
         LAYER m3 ;
         RECT  18.8 218.4 19.6 219.2 ;
         LAYER m3 ;
         RECT  181.3 306.1 181.9 306.7 ;
         LAYER m3 ;
         RECT  208.5 202.1 209.1 202.7 ;
         LAYER m3 ;
         RECT  181.3 326.9 181.9 327.5 ;
         LAYER m3 ;
         RECT  188.0 243.6 188.8 244.4 ;
         LAYER m3 ;
         RECT  208.5 222.9 209.1 223.5 ;
         LAYER m3 ;
         RECT  208.5 243.7 209.1 244.3 ;
         LAYER m3 ;
         RECT  144.7 285.6 145.5 286.4 ;
         LAYER m3 ;
         RECT  201.7 285.3 202.3 285.9 ;
         LAYER m3 ;
         RECT  181.3 243.7 181.9 244.3 ;
         LAYER m3 ;
         RECT  12.4 173.6 13.2 174.4 ;
         LAYER m3 ;
         RECT  181.3 347.7 181.9 348.3 ;
         LAYER m3 ;
         RECT  181.3 368.5 181.9 369.1 ;
         LAYER m3 ;
         RECT  6.0 218.4 6.8 219.2 ;
         LAYER m3 ;
         RECT  188.0 326.8 188.8 327.6 ;
         LAYER m3 ;
         RECT  118.7 202.4 119.5 203.2 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  205.1 280.3 205.7 280.9 ;
         LAYER m3 ;
         RECT  205.1 259.5 205.7 260.1 ;
         LAYER m3 ;
         RECT  198.3 259.5 198.9 260.1 ;
         LAYER m3 ;
         RECT  165.5 212.8 166.3 213.6 ;
         LAYER m3 ;
         RECT  184.7 186.3 185.3 186.9 ;
         LAYER m3 ;
         RECT  103.7 275.2 104.5 276.0 ;
         LAYER m3 ;
         RECT  184.6 363.4 185.4 364.2 ;
         LAYER m3 ;
         RECT  191.4 352.6 192.2 353.4 ;
         LAYER m3 ;
         RECT  184.6 290.2 185.4 291.0 ;
         LAYER m3 ;
         RECT  198.3 207.1 198.9 207.7 ;
         LAYER m3 ;
         RECT  184.6 207.0 185.4 207.8 ;
         LAYER m3 ;
         RECT  205.1 207.1 205.7 207.7 ;
         LAYER m3 ;
         RECT  184.7 280.3 185.3 280.9 ;
         LAYER m3 ;
         RECT  211.9 186.3 212.5 186.9 ;
         LAYER m3 ;
         RECT  103.7 233.6 104.5 234.4 ;
         LAYER m3 ;
         RECT  177.9 311.1 178.5 311.7 ;
         LAYER m3 ;
         RECT  205.1 269.5 205.7 270.1 ;
         LAYER m3 ;
         RECT  184.6 259.4 185.4 260.2 ;
         LAYER m3 ;
         RECT  191.5 186.3 192.1 186.9 ;
         LAYER m3 ;
         RECT  118.7 192.0 119.5 192.8 ;
         LAYER m3 ;
         RECT  165.5 358.4 166.3 359.2 ;
         LAYER m3 ;
         RECT  197.0 90.0 197.8 90.8 ;
         LAYER m3 ;
         RECT  191.4 321.8 192.2 322.6 ;
         LAYER m3 ;
         RECT  211.9 259.5 212.5 260.1 ;
         LAYER m3 ;
         RECT  184.6 238.6 185.4 239.4 ;
         LAYER m3 ;
         RECT  198.2 143.8 199.0 144.6 ;
         LAYER m3 ;
         RECT  211.9 342.7 212.5 343.3 ;
         LAYER m3 ;
         RECT  211.9 227.9 212.5 228.5 ;
         LAYER m3 ;
         RECT  177.9 259.5 178.5 260.1 ;
         LAYER m3 ;
         RECT  177.9 197.1 178.5 197.7 ;
         LAYER m3 ;
         RECT  144.7 358.4 145.5 359.2 ;
         LAYER m3 ;
         RECT  184.7 248.7 185.3 249.3 ;
         LAYER m3 ;
         RECT  103.7 212.8 104.5 213.6 ;
         LAYER m3 ;
         RECT  191.5 176.3 192.1 176.9 ;
         LAYER m3 ;
         RECT  191.5 248.7 192.1 249.3 ;
         LAYER m3 ;
         RECT  211.9 238.7 212.5 239.3 ;
         LAYER m3 ;
         RECT  205.1 217.9 205.7 218.5 ;
         LAYER m3 ;
         RECT  184.7 217.9 185.3 218.5 ;
         LAYER m3 ;
         RECT  191.4 311.0 192.2 311.8 ;
         LAYER m3 ;
         RECT  191.5 207.1 192.1 207.7 ;
         LAYER m3 ;
         RECT  191.5 197.1 192.1 197.7 ;
         LAYER m3 ;
         RECT  184.7 238.7 185.3 239.3 ;
         LAYER m3 ;
         RECT  144.7 296.0 145.5 296.8 ;
         LAYER m3 ;
         RECT  177.9 238.7 178.5 239.3 ;
         LAYER m3 ;
         RECT  6.0 252.0 6.8 252.8 ;
         LAYER m3 ;
         RECT  177.9 176.3 178.5 176.9 ;
         LAYER m3 ;
         RECT  191.5 259.5 192.1 260.1 ;
         LAYER m3 ;
         RECT  6.0 207.2 6.8 208.0 ;
         LAYER m3 ;
         RECT  211.9 290.3 212.5 290.9 ;
         LAYER m3 ;
         RECT  184.6 301.0 185.4 301.8 ;
         LAYER m3 ;
         RECT  205.1 331.9 205.7 332.5 ;
         LAYER m3 ;
         RECT  205.1 176.3 205.7 176.9 ;
         LAYER m3 ;
         RECT  191.5 269.5 192.1 270.1 ;
         LAYER m3 ;
         RECT  184.6 227.8 185.4 228.6 ;
         LAYER m3 ;
         RECT  191.4 363.4 192.2 364.2 ;
         LAYER m3 ;
         RECT  82.6 39.6 83.4 40.4 ;
         LAYER m3 ;
         RECT  191.5 321.9 192.1 322.5 ;
         LAYER m3 ;
         RECT  6.0 162.4 6.8 163.2 ;
         LAYER m3 ;
         RECT  18.8 162.4 19.6 163.2 ;
         LAYER m3 ;
         RECT  211.9 321.9 212.5 322.5 ;
         LAYER m3 ;
         RECT  191.4 248.6 192.2 249.4 ;
         LAYER m3 ;
         RECT  191.4 259.4 192.2 260.2 ;
         LAYER m3 ;
         RECT  205.1 363.5 205.7 364.1 ;
         LAYER m3 ;
         RECT  198.3 321.9 198.9 322.5 ;
         LAYER m3 ;
         RECT  82.6 119.6 83.4 120.4 ;
         LAYER m3 ;
         RECT  191.4 186.2 192.2 187.0 ;
         LAYER m3 ;
         RECT  177.9 227.9 178.5 228.5 ;
         LAYER m3 ;
         RECT  191.4 290.2 192.2 291.0 ;
         LAYER m3 ;
         RECT  184.7 311.1 185.3 311.7 ;
         LAYER m3 ;
         RECT  195.6 85.6 196.4 86.4 ;
         LAYER m3 ;
         RECT  177.9 248.7 178.5 249.3 ;
         LAYER m3 ;
         RECT  191.4 331.8 192.2 332.6 ;
         LAYER m3 ;
         RECT  198.3 331.9 198.9 332.5 ;
         LAYER m3 ;
         RECT  191.5 331.9 192.1 332.5 ;
         LAYER m3 ;
         RECT  184.6 248.6 185.4 249.4 ;
         LAYER m3 ;
         RECT  211.9 301.1 212.5 301.7 ;
         LAYER m3 ;
         RECT  205.1 186.3 205.7 186.9 ;
         LAYER m3 ;
         RECT  6.0 229.6 6.8 230.4 ;
         LAYER m3 ;
         RECT  198.3 176.3 198.9 176.9 ;
         LAYER m3 ;
         RECT  12.4 207.2 13.2 208.0 ;
         LAYER m3 ;
         RECT  144.7 316.8 145.5 317.6 ;
         LAYER m3 ;
         RECT  18.8 229.6 19.6 230.4 ;
         LAYER m3 ;
         RECT  198.3 269.5 198.9 270.1 ;
         LAYER m3 ;
         RECT  211.9 269.5 212.5 270.1 ;
         LAYER m3 ;
         RECT  118.7 233.6 119.5 234.4 ;
         LAYER m3 ;
         RECT  184.7 197.1 185.3 197.7 ;
         LAYER m3 ;
         RECT  118.7 254.4 119.5 255.2 ;
         LAYER m3 ;
         RECT  211.9 352.7 212.5 353.3 ;
         LAYER m3 ;
         RECT  198.3 197.1 198.9 197.7 ;
         LAYER m3 ;
         RECT  184.6 331.8 185.4 332.6 ;
         LAYER m3 ;
         RECT  165.5 192.0 166.3 192.8 ;
         LAYER m3 ;
         RECT  205.1 227.9 205.7 228.5 ;
         LAYER m3 ;
         RECT  211.9 197.1 212.5 197.7 ;
         LAYER m3 ;
         RECT  198.3 301.1 198.9 301.7 ;
         LAYER m3 ;
         RECT  191.4 342.6 192.2 343.4 ;
         LAYER m3 ;
         RECT  198.3 186.3 198.9 186.9 ;
         LAYER m3 ;
         RECT  118.7 212.8 119.5 213.6 ;
         LAYER m3 ;
         RECT  73.1 290.2 73.9 291.0 ;
         LAYER m3 ;
         RECT  202.4 85.6 203.2 86.4 ;
         LAYER m3 ;
         RECT  198.3 238.7 198.9 239.3 ;
         LAYER m3 ;
         RECT  210.5 45.4 211.3 46.2 ;
         LAYER m3 ;
         RECT  -0.4 39.6 0.4 40.4 ;
         LAYER m3 ;
         RECT  191.4 197.0 192.2 197.8 ;
         LAYER m3 ;
         RECT  205.1 352.7 205.7 353.3 ;
         LAYER m3 ;
         RECT  205.1 321.9 205.7 322.5 ;
         LAYER m3 ;
         RECT  191.5 217.9 192.1 218.5 ;
         LAYER m3 ;
         RECT  184.6 280.2 185.4 281.0 ;
         LAYER m3 ;
         RECT  194.2 104.6 195.0 105.4 ;
         LAYER m3 ;
         RECT  184.7 331.9 185.3 332.5 ;
         LAYER m3 ;
         RECT  184.6 269.4 185.4 270.2 ;
         LAYER m3 ;
         RECT  191.5 280.3 192.1 280.9 ;
         LAYER m3 ;
         RECT  198.3 311.1 198.9 311.7 ;
         LAYER m3 ;
         RECT  184.7 290.3 185.3 290.9 ;
         LAYER m3 ;
         RECT  191.4 238.6 192.2 239.4 ;
         LAYER m3 ;
         RECT  177.9 363.5 178.5 364.1 ;
         LAYER m3 ;
         RECT  184.6 311.0 185.4 311.8 ;
         LAYER m3 ;
         RECT  191.4 207.0 192.2 207.8 ;
         LAYER m3 ;
         RECT  198.3 363.5 198.9 364.1 ;
         LAYER m3 ;
         RECT  198.3 280.3 198.9 280.9 ;
         LAYER m3 ;
         RECT  73.1 330.2 73.9 331.0 ;
         LAYER m3 ;
         RECT  191.4 269.4 192.2 270.2 ;
         LAYER m3 ;
         RECT  211.9 363.5 212.5 364.1 ;
         LAYER m3 ;
         RECT  205.1 342.7 205.7 343.3 ;
         LAYER m3 ;
         RECT  177.9 186.3 178.5 186.9 ;
         LAYER m3 ;
         RECT  191.5 352.7 192.1 353.3 ;
         LAYER m3 ;
         RECT  18.8 207.2 19.6 208.0 ;
         LAYER m3 ;
         RECT  184.7 207.1 185.3 207.7 ;
         LAYER m3 ;
         RECT  82.6 -0.4 83.4 0.4 ;
         LAYER m3 ;
         RECT  191.5 227.9 192.1 228.5 ;
         LAYER m3 ;
         RECT  12.4 229.6 13.2 230.4 ;
         LAYER m3 ;
         RECT  12.4 162.4 13.2 163.2 ;
         LAYER m3 ;
         RECT  184.6 342.6 185.4 343.4 ;
         LAYER m3 ;
         RECT  211.9 248.7 212.5 249.3 ;
         LAYER m3 ;
         RECT  203.8 90.0 204.6 90.8 ;
         LAYER m3 ;
         RECT  6.0 184.8 6.8 185.6 ;
         LAYER m3 ;
         RECT  177.9 207.1 178.5 207.7 ;
         LAYER m3 ;
         RECT  177.9 342.7 178.5 343.3 ;
         LAYER m3 ;
         RECT  18.8 252.0 19.6 252.8 ;
         LAYER m3 ;
         RECT  198.3 217.9 198.9 218.5 ;
         LAYER m3 ;
         RECT  144.7 254.4 145.5 255.2 ;
         LAYER m3 ;
         RECT  184.6 176.2 185.4 177.0 ;
         LAYER m3 ;
         RECT  184.7 269.5 185.3 270.1 ;
         LAYER m3 ;
         RECT  177.9 280.3 178.5 280.9 ;
         LAYER m3 ;
         RECT  82.6 79.6 83.4 80.4 ;
         LAYER m3 ;
         RECT  191.5 238.7 192.1 239.3 ;
         LAYER m3 ;
         RECT  165.5 337.6 166.3 338.4 ;
         LAYER m3 ;
         RECT  205.1 248.7 205.7 249.3 ;
         LAYER m3 ;
         RECT  191.4 217.8 192.2 218.6 ;
         LAYER m3 ;
         RECT  211.9 207.1 212.5 207.7 ;
         LAYER m3 ;
         RECT  184.7 363.5 185.3 364.1 ;
         LAYER m3 ;
         RECT  144.7 275.2 145.5 276.0 ;
         LAYER m3 ;
         RECT  165.5 275.2 166.3 276.0 ;
         LAYER m3 ;
         RECT  211.9 176.3 212.5 176.9 ;
         LAYER m3 ;
         RECT  191.5 363.5 192.1 364.1 ;
         LAYER m3 ;
         RECT  198.3 248.7 198.9 249.3 ;
         LAYER m3 ;
         RECT  184.7 321.9 185.3 322.5 ;
         LAYER m3 ;
         RECT  191.4 280.2 192.2 281.0 ;
         LAYER m3 ;
         RECT  191.5 301.1 192.1 301.7 ;
         LAYER m3 ;
         RECT  165.5 296.0 166.3 296.8 ;
         LAYER m3 ;
         RECT  188.7 45.4 189.5 46.2 ;
         LAYER m3 ;
         RECT  103.7 192.0 104.5 192.8 ;
         LAYER m3 ;
         RECT  177.9 301.1 178.5 301.7 ;
         LAYER m3 ;
         RECT  205.0 143.8 205.8 144.6 ;
         LAYER m3 ;
         RECT  191.4 227.8 192.2 228.6 ;
         LAYER m3 ;
         RECT  205.1 238.7 205.7 239.3 ;
         LAYER m3 ;
         RECT  184.6 321.8 185.4 322.6 ;
         LAYER m3 ;
         RECT  144.7 212.8 145.5 213.6 ;
         LAYER m3 ;
         RECT  205.1 301.1 205.7 301.7 ;
         LAYER m3 ;
         RECT  177.9 217.9 178.5 218.5 ;
         LAYER m3 ;
         RECT  184.7 301.1 185.3 301.7 ;
         LAYER m3 ;
         RECT  73.1 370.2 73.9 371.0 ;
         LAYER m3 ;
         RECT  177.9 321.9 178.5 322.5 ;
         LAYER m3 ;
         RECT  12.4 184.8 13.2 185.6 ;
         LAYER m3 ;
         RECT  191.4 176.2 192.2 177.0 ;
         LAYER m3 ;
         RECT  184.6 197.0 185.4 197.8 ;
         LAYER m3 ;
         RECT  184.7 227.9 185.3 228.5 ;
         LAYER m3 ;
         RECT  198.3 352.7 198.9 353.3 ;
         LAYER m3 ;
         RECT  184.6 352.6 185.4 353.4 ;
         LAYER m3 ;
         RECT  184.7 352.7 185.3 353.3 ;
         LAYER m3 ;
         RECT  211.9 311.1 212.5 311.7 ;
         LAYER m3 ;
         RECT  144.7 192.0 145.5 192.8 ;
         LAYER m3 ;
         RECT  191.5 342.7 192.1 343.3 ;
         LAYER m3 ;
         RECT  201.0 104.6 201.8 105.4 ;
         LAYER m3 ;
         RECT  184.7 176.3 185.3 176.9 ;
         LAYER m3 ;
         RECT  118.7 275.2 119.5 276.0 ;
         LAYER m3 ;
         RECT  205.1 311.1 205.7 311.7 ;
         LAYER m3 ;
         RECT  184.6 186.2 185.4 187.0 ;
         LAYER m3 ;
         RECT  165.5 316.8 166.3 317.6 ;
         LAYER m3 ;
         RECT  177.9 269.5 178.5 270.1 ;
         LAYER m3 ;
         RECT  165.5 233.6 166.3 234.4 ;
         LAYER m3 ;
         RECT  165.5 254.4 166.3 255.2 ;
         LAYER m3 ;
         RECT  12.4 252.0 13.2 252.8 ;
         LAYER m3 ;
         RECT  184.7 259.5 185.3 260.1 ;
         LAYER m3 ;
         RECT  205.1 290.3 205.7 290.9 ;
         LAYER m3 ;
         RECT  184.7 342.7 185.3 343.3 ;
         LAYER m3 ;
         RECT  82.6 159.6 83.4 160.4 ;
         LAYER m3 ;
         RECT  211.9 331.9 212.5 332.5 ;
         LAYER m3 ;
         RECT  211.9 217.9 212.5 218.5 ;
         LAYER m3 ;
         RECT  191.5 290.3 192.1 290.9 ;
         LAYER m3 ;
         RECT  18.8 184.8 19.6 185.6 ;
         LAYER m3 ;
         RECT  211.9 280.3 212.5 280.9 ;
         LAYER m3 ;
         RECT  177.9 290.3 178.5 290.9 ;
         LAYER m3 ;
         RECT  177.9 331.9 178.5 332.5 ;
         LAYER m3 ;
         RECT  191.4 301.0 192.2 301.8 ;
         LAYER m3 ;
         RECT  198.3 342.7 198.9 343.3 ;
         LAYER m3 ;
         RECT  205.1 197.1 205.7 197.7 ;
         LAYER m3 ;
         RECT  103.7 254.4 104.5 255.2 ;
         LAYER m3 ;
         RECT  198.3 290.3 198.9 290.9 ;
         LAYER m3 ;
         RECT  144.7 233.6 145.5 234.4 ;
         LAYER m3 ;
         RECT  198.3 227.9 198.9 228.5 ;
         LAYER m3 ;
         RECT  191.5 311.1 192.1 311.7 ;
         LAYER m3 ;
         RECT  184.6 217.8 185.4 218.6 ;
         LAYER m3 ;
         RECT  144.7 337.6 145.5 338.4 ;
         LAYER m3 ;
         RECT  177.9 352.7 178.5 353.3 ;
         LAYER m3 ;
         RECT  -0.4 -0.4 0.4 0.4 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  191.4 202.0 199.0 202.8 ;
      RECT  198.2 200.4 199.0 202.0 ;
      RECT  196.4 196.8 197.2 197.2 ;
      RECT  193.0 192.8 194.6 193.6 ;
      RECT  196.4 198.0 197.2 200.4 ;
      RECT  191.4 194.2 199.0 195.0 ;
      RECT  195.2 195.0 196.0 195.2 ;
      RECT  194.0 200.4 195.0 201.2 ;
      RECT  191.4 195.6 192.2 199.8 ;
      RECT  194.0 199.8 194.8 200.4 ;
      RECT  191.4 200.4 192.2 202.0 ;
      RECT  196.0 197.2 197.2 198.0 ;
      RECT  195.8 192.8 197.4 193.6 ;
      RECT  196.4 196.0 197.4 196.8 ;
      RECT  196.2 200.4 197.2 201.2 ;
      RECT  193.8 196.0 194.8 196.8 ;
      RECT  194.0 196.8 194.8 199.0 ;
      RECT  194.0 199.0 195.6 199.8 ;
      RECT  198.2 195.6 199.0 199.8 ;
      RECT  191.4 202.8 199.0 202.0 ;
      RECT  198.2 204.4 199.0 202.8 ;
      RECT  196.4 208.0 197.2 207.6 ;
      RECT  193.0 212.0 194.6 211.2 ;
      RECT  196.4 206.8 197.2 204.4 ;
      RECT  191.4 210.6 199.0 209.8 ;
      RECT  195.2 209.8 196.0 209.6 ;
      RECT  194.0 204.4 195.0 203.6 ;
      RECT  191.4 209.2 192.2 205.0 ;
      RECT  194.0 205.0 194.8 204.4 ;
      RECT  191.4 204.4 192.2 202.8 ;
      RECT  196.0 207.6 197.2 206.8 ;
      RECT  195.8 212.0 197.4 211.2 ;
      RECT  196.4 208.8 197.4 208.0 ;
      RECT  196.2 204.4 197.2 203.6 ;
      RECT  193.8 208.8 194.8 208.0 ;
      RECT  194.0 208.0 194.8 205.8 ;
      RECT  194.0 205.8 195.6 205.0 ;
      RECT  198.2 209.2 199.0 205.0 ;
      RECT  191.4 222.8 199.0 223.6 ;
      RECT  198.2 221.2 199.0 222.8 ;
      RECT  196.4 217.6 197.2 218.0 ;
      RECT  193.0 213.6 194.6 214.4 ;
      RECT  196.4 218.8 197.2 221.2 ;
      RECT  191.4 215.0 199.0 215.8 ;
      RECT  195.2 215.8 196.0 216.0 ;
      RECT  194.0 221.2 195.0 222.0 ;
      RECT  191.4 216.4 192.2 220.6 ;
      RECT  194.0 220.6 194.8 221.2 ;
      RECT  191.4 221.2 192.2 222.8 ;
      RECT  196.0 218.0 197.2 218.8 ;
      RECT  195.8 213.6 197.4 214.4 ;
      RECT  196.4 216.8 197.4 217.6 ;
      RECT  196.2 221.2 197.2 222.0 ;
      RECT  193.8 216.8 194.8 217.6 ;
      RECT  194.0 217.6 194.8 219.8 ;
      RECT  194.0 219.8 195.6 220.6 ;
      RECT  198.2 216.4 199.0 220.6 ;
      RECT  191.4 223.6 199.0 222.8 ;
      RECT  198.2 225.2 199.0 223.6 ;
      RECT  196.4 228.8 197.2 228.4 ;
      RECT  193.0 232.8 194.6 232.0 ;
      RECT  196.4 227.6 197.2 225.2 ;
      RECT  191.4 231.4 199.0 230.6 ;
      RECT  195.2 230.6 196.0 230.4 ;
      RECT  194.0 225.2 195.0 224.4 ;
      RECT  191.4 230.0 192.2 225.8 ;
      RECT  194.0 225.8 194.8 225.2 ;
      RECT  191.4 225.2 192.2 223.6 ;
      RECT  196.0 228.4 197.2 227.6 ;
      RECT  195.8 232.8 197.4 232.0 ;
      RECT  196.4 229.6 197.4 228.8 ;
      RECT  196.2 225.2 197.2 224.4 ;
      RECT  193.8 229.6 194.8 228.8 ;
      RECT  194.0 228.8 194.8 226.6 ;
      RECT  194.0 226.6 195.6 225.8 ;
      RECT  198.2 230.0 199.0 225.8 ;
      RECT  191.4 243.6 199.0 244.4 ;
      RECT  198.2 242.0 199.0 243.6 ;
      RECT  196.4 238.4 197.2 238.8 ;
      RECT  193.0 234.4 194.6 235.2 ;
      RECT  196.4 239.6 197.2 242.0 ;
      RECT  191.4 235.8 199.0 236.6 ;
      RECT  195.2 236.6 196.0 236.8 ;
      RECT  194.0 242.0 195.0 242.8 ;
      RECT  191.4 237.2 192.2 241.4 ;
      RECT  194.0 241.4 194.8 242.0 ;
      RECT  191.4 242.0 192.2 243.6 ;
      RECT  196.0 238.8 197.2 239.6 ;
      RECT  195.8 234.4 197.4 235.2 ;
      RECT  196.4 237.6 197.4 238.4 ;
      RECT  196.2 242.0 197.2 242.8 ;
      RECT  193.8 237.6 194.8 238.4 ;
      RECT  194.0 238.4 194.8 240.6 ;
      RECT  194.0 240.6 195.6 241.4 ;
      RECT  198.2 237.2 199.0 241.4 ;
      RECT  191.4 244.4 199.0 243.6 ;
      RECT  198.2 246.0 199.0 244.4 ;
      RECT  196.4 249.6 197.2 249.2 ;
      RECT  193.0 253.6 194.6 252.8 ;
      RECT  196.4 248.4 197.2 246.0 ;
      RECT  191.4 252.2 199.0 251.4 ;
      RECT  195.2 251.4 196.0 251.2 ;
      RECT  194.0 246.0 195.0 245.2 ;
      RECT  191.4 250.8 192.2 246.6 ;
      RECT  194.0 246.6 194.8 246.0 ;
      RECT  191.4 246.0 192.2 244.4 ;
      RECT  196.0 249.2 197.2 248.4 ;
      RECT  195.8 253.6 197.4 252.8 ;
      RECT  196.4 250.4 197.4 249.6 ;
      RECT  196.2 246.0 197.2 245.2 ;
      RECT  193.8 250.4 194.8 249.6 ;
      RECT  194.0 249.6 194.8 247.4 ;
      RECT  194.0 247.4 195.6 246.6 ;
      RECT  198.2 250.8 199.0 246.6 ;
      RECT  191.4 264.4 199.0 265.2 ;
      RECT  198.2 262.8 199.0 264.4 ;
      RECT  196.4 259.2 197.2 259.6 ;
      RECT  193.0 255.2 194.6 256.0 ;
      RECT  196.4 260.4 197.2 262.8 ;
      RECT  191.4 256.6 199.0 257.4 ;
      RECT  195.2 257.4 196.0 257.6 ;
      RECT  194.0 262.8 195.0 263.6 ;
      RECT  191.4 258.0 192.2 262.2 ;
      RECT  194.0 262.2 194.8 262.8 ;
      RECT  191.4 262.8 192.2 264.4 ;
      RECT  196.0 259.6 197.2 260.4 ;
      RECT  195.8 255.2 197.4 256.0 ;
      RECT  196.4 258.4 197.4 259.2 ;
      RECT  196.2 262.8 197.2 263.6 ;
      RECT  193.8 258.4 194.8 259.2 ;
      RECT  194.0 259.2 194.8 261.4 ;
      RECT  194.0 261.4 195.6 262.2 ;
      RECT  198.2 258.0 199.0 262.2 ;
      RECT  191.4 265.2 199.0 264.4 ;
      RECT  198.2 266.8 199.0 265.2 ;
      RECT  196.4 270.4 197.2 270.0 ;
      RECT  193.0 274.4 194.6 273.6 ;
      RECT  196.4 269.2 197.2 266.8 ;
      RECT  191.4 273.0 199.0 272.2 ;
      RECT  195.2 272.2 196.0 272.0 ;
      RECT  194.0 266.8 195.0 266.0 ;
      RECT  191.4 271.6 192.2 267.4 ;
      RECT  194.0 267.4 194.8 266.8 ;
      RECT  191.4 266.8 192.2 265.2 ;
      RECT  196.0 270.0 197.2 269.2 ;
      RECT  195.8 274.4 197.4 273.6 ;
      RECT  196.4 271.2 197.4 270.4 ;
      RECT  196.2 266.8 197.2 266.0 ;
      RECT  193.8 271.2 194.8 270.4 ;
      RECT  194.0 270.4 194.8 268.2 ;
      RECT  194.0 268.2 195.6 267.4 ;
      RECT  198.2 271.6 199.0 267.4 ;
      RECT  191.4 285.2 199.0 286.0 ;
      RECT  198.2 283.6 199.0 285.2 ;
      RECT  196.4 280.0 197.2 280.4 ;
      RECT  193.0 276.0 194.6 276.8 ;
      RECT  196.4 281.2 197.2 283.6 ;
      RECT  191.4 277.4 199.0 278.2 ;
      RECT  195.2 278.2 196.0 278.4 ;
      RECT  194.0 283.6 195.0 284.4 ;
      RECT  191.4 278.8 192.2 283.0 ;
      RECT  194.0 283.0 194.8 283.6 ;
      RECT  191.4 283.6 192.2 285.2 ;
      RECT  196.0 280.4 197.2 281.2 ;
      RECT  195.8 276.0 197.4 276.8 ;
      RECT  196.4 279.2 197.4 280.0 ;
      RECT  196.2 283.6 197.2 284.4 ;
      RECT  193.8 279.2 194.8 280.0 ;
      RECT  194.0 280.0 194.8 282.2 ;
      RECT  194.0 282.2 195.6 283.0 ;
      RECT  198.2 278.8 199.0 283.0 ;
      RECT  191.4 286.0 199.0 285.2 ;
      RECT  198.2 287.6 199.0 286.0 ;
      RECT  196.4 291.2 197.2 290.8 ;
      RECT  193.0 295.2 194.6 294.4 ;
      RECT  196.4 290.0 197.2 287.6 ;
      RECT  191.4 293.8 199.0 293.0 ;
      RECT  195.2 293.0 196.0 292.8 ;
      RECT  194.0 287.6 195.0 286.8 ;
      RECT  191.4 292.4 192.2 288.2 ;
      RECT  194.0 288.2 194.8 287.6 ;
      RECT  191.4 287.6 192.2 286.0 ;
      RECT  196.0 290.8 197.2 290.0 ;
      RECT  195.8 295.2 197.4 294.4 ;
      RECT  196.4 292.0 197.4 291.2 ;
      RECT  196.2 287.6 197.2 286.8 ;
      RECT  193.8 292.0 194.8 291.2 ;
      RECT  194.0 291.2 194.8 289.0 ;
      RECT  194.0 289.0 195.6 288.2 ;
      RECT  198.2 292.4 199.0 288.2 ;
      RECT  191.4 306.0 199.0 306.8 ;
      RECT  198.2 304.4 199.0 306.0 ;
      RECT  196.4 300.8 197.2 301.2 ;
      RECT  193.0 296.8 194.6 297.6 ;
      RECT  196.4 302.0 197.2 304.4 ;
      RECT  191.4 298.2 199.0 299.0 ;
      RECT  195.2 299.0 196.0 299.2 ;
      RECT  194.0 304.4 195.0 305.2 ;
      RECT  191.4 299.6 192.2 303.8 ;
      RECT  194.0 303.8 194.8 304.4 ;
      RECT  191.4 304.4 192.2 306.0 ;
      RECT  196.0 301.2 197.2 302.0 ;
      RECT  195.8 296.8 197.4 297.6 ;
      RECT  196.4 300.0 197.4 300.8 ;
      RECT  196.2 304.4 197.2 305.2 ;
      RECT  193.8 300.0 194.8 300.8 ;
      RECT  194.0 300.8 194.8 303.0 ;
      RECT  194.0 303.0 195.6 303.8 ;
      RECT  198.2 299.6 199.0 303.8 ;
      RECT  191.4 306.8 199.0 306.0 ;
      RECT  198.2 308.4 199.0 306.8 ;
      RECT  196.4 312.0 197.2 311.6 ;
      RECT  193.0 316.0 194.6 315.2 ;
      RECT  196.4 310.8 197.2 308.4 ;
      RECT  191.4 314.6 199.0 313.8 ;
      RECT  195.2 313.8 196.0 313.6 ;
      RECT  194.0 308.4 195.0 307.6 ;
      RECT  191.4 313.2 192.2 309.0 ;
      RECT  194.0 309.0 194.8 308.4 ;
      RECT  191.4 308.4 192.2 306.8 ;
      RECT  196.0 311.6 197.2 310.8 ;
      RECT  195.8 316.0 197.4 315.2 ;
      RECT  196.4 312.8 197.4 312.0 ;
      RECT  196.2 308.4 197.2 307.6 ;
      RECT  193.8 312.8 194.8 312.0 ;
      RECT  194.0 312.0 194.8 309.8 ;
      RECT  194.0 309.8 195.6 309.0 ;
      RECT  198.2 313.2 199.0 309.0 ;
      RECT  191.4 326.8 199.0 327.6 ;
      RECT  198.2 325.2 199.0 326.8 ;
      RECT  196.4 321.6 197.2 322.0 ;
      RECT  193.0 317.6 194.6 318.4 ;
      RECT  196.4 322.8 197.2 325.2 ;
      RECT  191.4 319.0 199.0 319.8 ;
      RECT  195.2 319.8 196.0 320.0 ;
      RECT  194.0 325.2 195.0 326.0 ;
      RECT  191.4 320.4 192.2 324.6 ;
      RECT  194.0 324.6 194.8 325.2 ;
      RECT  191.4 325.2 192.2 326.8 ;
      RECT  196.0 322.0 197.2 322.8 ;
      RECT  195.8 317.6 197.4 318.4 ;
      RECT  196.4 320.8 197.4 321.6 ;
      RECT  196.2 325.2 197.2 326.0 ;
      RECT  193.8 320.8 194.8 321.6 ;
      RECT  194.0 321.6 194.8 323.8 ;
      RECT  194.0 323.8 195.6 324.6 ;
      RECT  198.2 320.4 199.0 324.6 ;
      RECT  191.4 327.6 199.0 326.8 ;
      RECT  198.2 329.2 199.0 327.6 ;
      RECT  196.4 332.8 197.2 332.4 ;
      RECT  193.0 336.8 194.6 336.0 ;
      RECT  196.4 331.6 197.2 329.2 ;
      RECT  191.4 335.4 199.0 334.6 ;
      RECT  195.2 334.6 196.0 334.4 ;
      RECT  194.0 329.2 195.0 328.4 ;
      RECT  191.4 334.0 192.2 329.8 ;
      RECT  194.0 329.8 194.8 329.2 ;
      RECT  191.4 329.2 192.2 327.6 ;
      RECT  196.0 332.4 197.2 331.6 ;
      RECT  195.8 336.8 197.4 336.0 ;
      RECT  196.4 333.6 197.4 332.8 ;
      RECT  196.2 329.2 197.2 328.4 ;
      RECT  193.8 333.6 194.8 332.8 ;
      RECT  194.0 332.8 194.8 330.6 ;
      RECT  194.0 330.6 195.6 329.8 ;
      RECT  198.2 334.0 199.0 329.8 ;
      RECT  191.4 347.6 199.0 348.4 ;
      RECT  198.2 346.0 199.0 347.6 ;
      RECT  196.4 342.4 197.2 342.8 ;
      RECT  193.0 338.4 194.6 339.2 ;
      RECT  196.4 343.6 197.2 346.0 ;
      RECT  191.4 339.8 199.0 340.6 ;
      RECT  195.2 340.6 196.0 340.8 ;
      RECT  194.0 346.0 195.0 346.8 ;
      RECT  191.4 341.2 192.2 345.4 ;
      RECT  194.0 345.4 194.8 346.0 ;
      RECT  191.4 346.0 192.2 347.6 ;
      RECT  196.0 342.8 197.2 343.6 ;
      RECT  195.8 338.4 197.4 339.2 ;
      RECT  196.4 341.6 197.4 342.4 ;
      RECT  196.2 346.0 197.2 346.8 ;
      RECT  193.8 341.6 194.8 342.4 ;
      RECT  194.0 342.4 194.8 344.6 ;
      RECT  194.0 344.6 195.6 345.4 ;
      RECT  198.2 341.2 199.0 345.4 ;
      RECT  191.4 348.4 199.0 347.6 ;
      RECT  198.2 350.0 199.0 348.4 ;
      RECT  196.4 353.6 197.2 353.2 ;
      RECT  193.0 357.6 194.6 356.8 ;
      RECT  196.4 352.4 197.2 350.0 ;
      RECT  191.4 356.2 199.0 355.4 ;
      RECT  195.2 355.4 196.0 355.2 ;
      RECT  194.0 350.0 195.0 349.2 ;
      RECT  191.4 354.8 192.2 350.6 ;
      RECT  194.0 350.6 194.8 350.0 ;
      RECT  191.4 350.0 192.2 348.4 ;
      RECT  196.0 353.2 197.2 352.4 ;
      RECT  195.8 357.6 197.4 356.8 ;
      RECT  196.4 354.4 197.4 353.6 ;
      RECT  196.2 350.0 197.2 349.2 ;
      RECT  193.8 354.4 194.8 353.6 ;
      RECT  194.0 353.6 194.8 351.4 ;
      RECT  194.0 351.4 195.6 350.6 ;
      RECT  198.2 354.8 199.0 350.6 ;
      RECT  198.2 202.0 205.8 202.8 ;
      RECT  205.0 200.4 205.8 202.0 ;
      RECT  203.2 196.8 204.0 197.2 ;
      RECT  199.8 192.8 201.4 193.6 ;
      RECT  203.2 198.0 204.0 200.4 ;
      RECT  198.2 194.2 205.8 195.0 ;
      RECT  202.0 195.0 202.8 195.2 ;
      RECT  200.8 200.4 201.8 201.2 ;
      RECT  198.2 195.6 199.0 199.8 ;
      RECT  200.8 199.8 201.6 200.4 ;
      RECT  198.2 200.4 199.0 202.0 ;
      RECT  202.8 197.2 204.0 198.0 ;
      RECT  202.6 192.8 204.2 193.6 ;
      RECT  203.2 196.0 204.2 196.8 ;
      RECT  203.0 200.4 204.0 201.2 ;
      RECT  200.6 196.0 201.6 196.8 ;
      RECT  200.8 196.8 201.6 199.0 ;
      RECT  200.8 199.0 202.4 199.8 ;
      RECT  205.0 195.6 205.8 199.8 ;
      RECT  198.2 202.8 205.8 202.0 ;
      RECT  205.0 204.4 205.8 202.8 ;
      RECT  203.2 208.0 204.0 207.6 ;
      RECT  199.8 212.0 201.4 211.2 ;
      RECT  203.2 206.8 204.0 204.4 ;
      RECT  198.2 210.6 205.8 209.8 ;
      RECT  202.0 209.8 202.8 209.6 ;
      RECT  200.8 204.4 201.8 203.6 ;
      RECT  198.2 209.2 199.0 205.0 ;
      RECT  200.8 205.0 201.6 204.4 ;
      RECT  198.2 204.4 199.0 202.8 ;
      RECT  202.8 207.6 204.0 206.8 ;
      RECT  202.6 212.0 204.2 211.2 ;
      RECT  203.2 208.8 204.2 208.0 ;
      RECT  203.0 204.4 204.0 203.6 ;
      RECT  200.6 208.8 201.6 208.0 ;
      RECT  200.8 208.0 201.6 205.8 ;
      RECT  200.8 205.8 202.4 205.0 ;
      RECT  205.0 209.2 205.8 205.0 ;
      RECT  198.2 222.8 205.8 223.6 ;
      RECT  205.0 221.2 205.8 222.8 ;
      RECT  203.2 217.6 204.0 218.0 ;
      RECT  199.8 213.6 201.4 214.4 ;
      RECT  203.2 218.8 204.0 221.2 ;
      RECT  198.2 215.0 205.8 215.8 ;
      RECT  202.0 215.8 202.8 216.0 ;
      RECT  200.8 221.2 201.8 222.0 ;
      RECT  198.2 216.4 199.0 220.6 ;
      RECT  200.8 220.6 201.6 221.2 ;
      RECT  198.2 221.2 199.0 222.8 ;
      RECT  202.8 218.0 204.0 218.8 ;
      RECT  202.6 213.6 204.2 214.4 ;
      RECT  203.2 216.8 204.2 217.6 ;
      RECT  203.0 221.2 204.0 222.0 ;
      RECT  200.6 216.8 201.6 217.6 ;
      RECT  200.8 217.6 201.6 219.8 ;
      RECT  200.8 219.8 202.4 220.6 ;
      RECT  205.0 216.4 205.8 220.6 ;
      RECT  198.2 223.6 205.8 222.8 ;
      RECT  205.0 225.2 205.8 223.6 ;
      RECT  203.2 228.8 204.0 228.4 ;
      RECT  199.8 232.8 201.4 232.0 ;
      RECT  203.2 227.6 204.0 225.2 ;
      RECT  198.2 231.4 205.8 230.6 ;
      RECT  202.0 230.6 202.8 230.4 ;
      RECT  200.8 225.2 201.8 224.4 ;
      RECT  198.2 230.0 199.0 225.8 ;
      RECT  200.8 225.8 201.6 225.2 ;
      RECT  198.2 225.2 199.0 223.6 ;
      RECT  202.8 228.4 204.0 227.6 ;
      RECT  202.6 232.8 204.2 232.0 ;
      RECT  203.2 229.6 204.2 228.8 ;
      RECT  203.0 225.2 204.0 224.4 ;
      RECT  200.6 229.6 201.6 228.8 ;
      RECT  200.8 228.8 201.6 226.6 ;
      RECT  200.8 226.6 202.4 225.8 ;
      RECT  205.0 230.0 205.8 225.8 ;
      RECT  198.2 243.6 205.8 244.4 ;
      RECT  205.0 242.0 205.8 243.6 ;
      RECT  203.2 238.4 204.0 238.8 ;
      RECT  199.8 234.4 201.4 235.2 ;
      RECT  203.2 239.6 204.0 242.0 ;
      RECT  198.2 235.8 205.8 236.6 ;
      RECT  202.0 236.6 202.8 236.8 ;
      RECT  200.8 242.0 201.8 242.8 ;
      RECT  198.2 237.2 199.0 241.4 ;
      RECT  200.8 241.4 201.6 242.0 ;
      RECT  198.2 242.0 199.0 243.6 ;
      RECT  202.8 238.8 204.0 239.6 ;
      RECT  202.6 234.4 204.2 235.2 ;
      RECT  203.2 237.6 204.2 238.4 ;
      RECT  203.0 242.0 204.0 242.8 ;
      RECT  200.6 237.6 201.6 238.4 ;
      RECT  200.8 238.4 201.6 240.6 ;
      RECT  200.8 240.6 202.4 241.4 ;
      RECT  205.0 237.2 205.8 241.4 ;
      RECT  198.2 244.4 205.8 243.6 ;
      RECT  205.0 246.0 205.8 244.4 ;
      RECT  203.2 249.6 204.0 249.2 ;
      RECT  199.8 253.6 201.4 252.8 ;
      RECT  203.2 248.4 204.0 246.0 ;
      RECT  198.2 252.2 205.8 251.4 ;
      RECT  202.0 251.4 202.8 251.2 ;
      RECT  200.8 246.0 201.8 245.2 ;
      RECT  198.2 250.8 199.0 246.6 ;
      RECT  200.8 246.6 201.6 246.0 ;
      RECT  198.2 246.0 199.0 244.4 ;
      RECT  202.8 249.2 204.0 248.4 ;
      RECT  202.6 253.6 204.2 252.8 ;
      RECT  203.2 250.4 204.2 249.6 ;
      RECT  203.0 246.0 204.0 245.2 ;
      RECT  200.6 250.4 201.6 249.6 ;
      RECT  200.8 249.6 201.6 247.4 ;
      RECT  200.8 247.4 202.4 246.6 ;
      RECT  205.0 250.8 205.8 246.6 ;
      RECT  198.2 264.4 205.8 265.2 ;
      RECT  205.0 262.8 205.8 264.4 ;
      RECT  203.2 259.2 204.0 259.6 ;
      RECT  199.8 255.2 201.4 256.0 ;
      RECT  203.2 260.4 204.0 262.8 ;
      RECT  198.2 256.6 205.8 257.4 ;
      RECT  202.0 257.4 202.8 257.6 ;
      RECT  200.8 262.8 201.8 263.6 ;
      RECT  198.2 258.0 199.0 262.2 ;
      RECT  200.8 262.2 201.6 262.8 ;
      RECT  198.2 262.8 199.0 264.4 ;
      RECT  202.8 259.6 204.0 260.4 ;
      RECT  202.6 255.2 204.2 256.0 ;
      RECT  203.2 258.4 204.2 259.2 ;
      RECT  203.0 262.8 204.0 263.6 ;
      RECT  200.6 258.4 201.6 259.2 ;
      RECT  200.8 259.2 201.6 261.4 ;
      RECT  200.8 261.4 202.4 262.2 ;
      RECT  205.0 258.0 205.8 262.2 ;
      RECT  198.2 265.2 205.8 264.4 ;
      RECT  205.0 266.8 205.8 265.2 ;
      RECT  203.2 270.4 204.0 270.0 ;
      RECT  199.8 274.4 201.4 273.6 ;
      RECT  203.2 269.2 204.0 266.8 ;
      RECT  198.2 273.0 205.8 272.2 ;
      RECT  202.0 272.2 202.8 272.0 ;
      RECT  200.8 266.8 201.8 266.0 ;
      RECT  198.2 271.6 199.0 267.4 ;
      RECT  200.8 267.4 201.6 266.8 ;
      RECT  198.2 266.8 199.0 265.2 ;
      RECT  202.8 270.0 204.0 269.2 ;
      RECT  202.6 274.4 204.2 273.6 ;
      RECT  203.2 271.2 204.2 270.4 ;
      RECT  203.0 266.8 204.0 266.0 ;
      RECT  200.6 271.2 201.6 270.4 ;
      RECT  200.8 270.4 201.6 268.2 ;
      RECT  200.8 268.2 202.4 267.4 ;
      RECT  205.0 271.6 205.8 267.4 ;
      RECT  198.2 285.2 205.8 286.0 ;
      RECT  205.0 283.6 205.8 285.2 ;
      RECT  203.2 280.0 204.0 280.4 ;
      RECT  199.8 276.0 201.4 276.8 ;
      RECT  203.2 281.2 204.0 283.6 ;
      RECT  198.2 277.4 205.8 278.2 ;
      RECT  202.0 278.2 202.8 278.4 ;
      RECT  200.8 283.6 201.8 284.4 ;
      RECT  198.2 278.8 199.0 283.0 ;
      RECT  200.8 283.0 201.6 283.6 ;
      RECT  198.2 283.6 199.0 285.2 ;
      RECT  202.8 280.4 204.0 281.2 ;
      RECT  202.6 276.0 204.2 276.8 ;
      RECT  203.2 279.2 204.2 280.0 ;
      RECT  203.0 283.6 204.0 284.4 ;
      RECT  200.6 279.2 201.6 280.0 ;
      RECT  200.8 280.0 201.6 282.2 ;
      RECT  200.8 282.2 202.4 283.0 ;
      RECT  205.0 278.8 205.8 283.0 ;
      RECT  198.2 286.0 205.8 285.2 ;
      RECT  205.0 287.6 205.8 286.0 ;
      RECT  203.2 291.2 204.0 290.8 ;
      RECT  199.8 295.2 201.4 294.4 ;
      RECT  203.2 290.0 204.0 287.6 ;
      RECT  198.2 293.8 205.8 293.0 ;
      RECT  202.0 293.0 202.8 292.8 ;
      RECT  200.8 287.6 201.8 286.8 ;
      RECT  198.2 292.4 199.0 288.2 ;
      RECT  200.8 288.2 201.6 287.6 ;
      RECT  198.2 287.6 199.0 286.0 ;
      RECT  202.8 290.8 204.0 290.0 ;
      RECT  202.6 295.2 204.2 294.4 ;
      RECT  203.2 292.0 204.2 291.2 ;
      RECT  203.0 287.6 204.0 286.8 ;
      RECT  200.6 292.0 201.6 291.2 ;
      RECT  200.8 291.2 201.6 289.0 ;
      RECT  200.8 289.0 202.4 288.2 ;
      RECT  205.0 292.4 205.8 288.2 ;
      RECT  198.2 306.0 205.8 306.8 ;
      RECT  205.0 304.4 205.8 306.0 ;
      RECT  203.2 300.8 204.0 301.2 ;
      RECT  199.8 296.8 201.4 297.6 ;
      RECT  203.2 302.0 204.0 304.4 ;
      RECT  198.2 298.2 205.8 299.0 ;
      RECT  202.0 299.0 202.8 299.2 ;
      RECT  200.8 304.4 201.8 305.2 ;
      RECT  198.2 299.6 199.0 303.8 ;
      RECT  200.8 303.8 201.6 304.4 ;
      RECT  198.2 304.4 199.0 306.0 ;
      RECT  202.8 301.2 204.0 302.0 ;
      RECT  202.6 296.8 204.2 297.6 ;
      RECT  203.2 300.0 204.2 300.8 ;
      RECT  203.0 304.4 204.0 305.2 ;
      RECT  200.6 300.0 201.6 300.8 ;
      RECT  200.8 300.8 201.6 303.0 ;
      RECT  200.8 303.0 202.4 303.8 ;
      RECT  205.0 299.6 205.8 303.8 ;
      RECT  198.2 306.8 205.8 306.0 ;
      RECT  205.0 308.4 205.8 306.8 ;
      RECT  203.2 312.0 204.0 311.6 ;
      RECT  199.8 316.0 201.4 315.2 ;
      RECT  203.2 310.8 204.0 308.4 ;
      RECT  198.2 314.6 205.8 313.8 ;
      RECT  202.0 313.8 202.8 313.6 ;
      RECT  200.8 308.4 201.8 307.6 ;
      RECT  198.2 313.2 199.0 309.0 ;
      RECT  200.8 309.0 201.6 308.4 ;
      RECT  198.2 308.4 199.0 306.8 ;
      RECT  202.8 311.6 204.0 310.8 ;
      RECT  202.6 316.0 204.2 315.2 ;
      RECT  203.2 312.8 204.2 312.0 ;
      RECT  203.0 308.4 204.0 307.6 ;
      RECT  200.6 312.8 201.6 312.0 ;
      RECT  200.8 312.0 201.6 309.8 ;
      RECT  200.8 309.8 202.4 309.0 ;
      RECT  205.0 313.2 205.8 309.0 ;
      RECT  198.2 326.8 205.8 327.6 ;
      RECT  205.0 325.2 205.8 326.8 ;
      RECT  203.2 321.6 204.0 322.0 ;
      RECT  199.8 317.6 201.4 318.4 ;
      RECT  203.2 322.8 204.0 325.2 ;
      RECT  198.2 319.0 205.8 319.8 ;
      RECT  202.0 319.8 202.8 320.0 ;
      RECT  200.8 325.2 201.8 326.0 ;
      RECT  198.2 320.4 199.0 324.6 ;
      RECT  200.8 324.6 201.6 325.2 ;
      RECT  198.2 325.2 199.0 326.8 ;
      RECT  202.8 322.0 204.0 322.8 ;
      RECT  202.6 317.6 204.2 318.4 ;
      RECT  203.2 320.8 204.2 321.6 ;
      RECT  203.0 325.2 204.0 326.0 ;
      RECT  200.6 320.8 201.6 321.6 ;
      RECT  200.8 321.6 201.6 323.8 ;
      RECT  200.8 323.8 202.4 324.6 ;
      RECT  205.0 320.4 205.8 324.6 ;
      RECT  198.2 327.6 205.8 326.8 ;
      RECT  205.0 329.2 205.8 327.6 ;
      RECT  203.2 332.8 204.0 332.4 ;
      RECT  199.8 336.8 201.4 336.0 ;
      RECT  203.2 331.6 204.0 329.2 ;
      RECT  198.2 335.4 205.8 334.6 ;
      RECT  202.0 334.6 202.8 334.4 ;
      RECT  200.8 329.2 201.8 328.4 ;
      RECT  198.2 334.0 199.0 329.8 ;
      RECT  200.8 329.8 201.6 329.2 ;
      RECT  198.2 329.2 199.0 327.6 ;
      RECT  202.8 332.4 204.0 331.6 ;
      RECT  202.6 336.8 204.2 336.0 ;
      RECT  203.2 333.6 204.2 332.8 ;
      RECT  203.0 329.2 204.0 328.4 ;
      RECT  200.6 333.6 201.6 332.8 ;
      RECT  200.8 332.8 201.6 330.6 ;
      RECT  200.8 330.6 202.4 329.8 ;
      RECT  205.0 334.0 205.8 329.8 ;
      RECT  198.2 347.6 205.8 348.4 ;
      RECT  205.0 346.0 205.8 347.6 ;
      RECT  203.2 342.4 204.0 342.8 ;
      RECT  199.8 338.4 201.4 339.2 ;
      RECT  203.2 343.6 204.0 346.0 ;
      RECT  198.2 339.8 205.8 340.6 ;
      RECT  202.0 340.6 202.8 340.8 ;
      RECT  200.8 346.0 201.8 346.8 ;
      RECT  198.2 341.2 199.0 345.4 ;
      RECT  200.8 345.4 201.6 346.0 ;
      RECT  198.2 346.0 199.0 347.6 ;
      RECT  202.8 342.8 204.0 343.6 ;
      RECT  202.6 338.4 204.2 339.2 ;
      RECT  203.2 341.6 204.2 342.4 ;
      RECT  203.0 346.0 204.0 346.8 ;
      RECT  200.6 341.6 201.6 342.4 ;
      RECT  200.8 342.4 201.6 344.6 ;
      RECT  200.8 344.6 202.4 345.4 ;
      RECT  205.0 341.2 205.8 345.4 ;
      RECT  198.2 348.4 205.8 347.6 ;
      RECT  205.0 350.0 205.8 348.4 ;
      RECT  203.2 353.6 204.0 353.2 ;
      RECT  199.8 357.6 201.4 356.8 ;
      RECT  203.2 352.4 204.0 350.0 ;
      RECT  198.2 356.2 205.8 355.4 ;
      RECT  202.0 355.4 202.8 355.2 ;
      RECT  200.8 350.0 201.8 349.2 ;
      RECT  198.2 354.8 199.0 350.6 ;
      RECT  200.8 350.6 201.6 350.0 ;
      RECT  198.2 350.0 199.0 348.4 ;
      RECT  202.8 353.2 204.0 352.4 ;
      RECT  202.6 357.6 204.2 356.8 ;
      RECT  203.2 354.4 204.2 353.6 ;
      RECT  203.0 350.0 204.0 349.2 ;
      RECT  200.6 354.4 201.6 353.6 ;
      RECT  200.8 353.6 201.6 351.4 ;
      RECT  200.8 351.4 202.4 350.6 ;
      RECT  205.0 354.8 205.8 350.6 ;
      RECT  191.8 194.2 205.4 195.0 ;
      RECT  191.8 209.8 205.4 210.6 ;
      RECT  191.8 215.0 205.4 215.8 ;
      RECT  191.8 230.6 205.4 231.4 ;
      RECT  191.8 235.8 205.4 236.6 ;
      RECT  191.8 251.4 205.4 252.2 ;
      RECT  191.8 256.6 205.4 257.4 ;
      RECT  191.8 272.2 205.4 273.0 ;
      RECT  191.8 277.4 205.4 278.2 ;
      RECT  191.8 293.0 205.4 293.8 ;
      RECT  191.8 298.2 205.4 299.0 ;
      RECT  191.8 313.8 205.4 314.6 ;
      RECT  191.8 319.0 205.4 319.8 ;
      RECT  191.8 334.6 205.4 335.4 ;
      RECT  191.8 339.8 205.4 340.6 ;
      RECT  191.8 355.4 205.4 356.2 ;
      RECT  184.6 181.2 192.2 182.0 ;
      RECT  191.4 179.6 192.2 181.2 ;
      RECT  189.6 176.0 190.4 176.4 ;
      RECT  189.6 177.2 190.4 179.6 ;
      RECT  184.6 173.4 192.2 174.2 ;
      RECT  189.8 172.0 190.6 172.8 ;
      RECT  188.4 174.2 189.2 174.4 ;
      RECT  187.2 179.6 188.2 180.4 ;
      RECT  184.6 174.8 185.4 179.0 ;
      RECT  187.2 179.0 188.0 179.6 ;
      RECT  184.6 179.6 185.4 181.2 ;
      RECT  189.2 176.4 190.4 177.2 ;
      RECT  189.6 175.2 190.6 176.0 ;
      RECT  189.4 179.6 190.4 180.4 ;
      RECT  187.0 175.2 188.0 176.0 ;
      RECT  187.2 176.0 188.0 178.2 ;
      RECT  187.2 178.2 188.8 179.0 ;
      RECT  187.0 172.0 187.8 172.8 ;
      RECT  191.4 174.8 192.2 179.0 ;
      RECT  184.6 182.0 192.2 181.2 ;
      RECT  191.4 183.6 192.2 182.0 ;
      RECT  189.6 187.2 190.4 186.8 ;
      RECT  186.2 191.2 187.8 190.4 ;
      RECT  189.6 186.0 190.4 183.6 ;
      RECT  184.6 189.8 192.2 189.0 ;
      RECT  189.4 182.8 190.2 182.0 ;
      RECT  188.4 189.0 189.2 188.8 ;
      RECT  187.2 183.6 188.2 182.8 ;
      RECT  184.6 188.4 185.4 184.2 ;
      RECT  187.2 184.2 188.0 183.6 ;
      RECT  184.6 183.6 185.4 182.0 ;
      RECT  189.2 186.8 190.4 186.0 ;
      RECT  189.0 191.2 190.6 190.4 ;
      RECT  189.6 188.0 190.6 187.2 ;
      RECT  189.4 183.6 190.4 182.8 ;
      RECT  187.0 188.0 188.0 187.2 ;
      RECT  187.2 187.2 188.0 185.0 ;
      RECT  187.2 185.0 188.8 184.2 ;
      RECT  191.4 188.4 192.2 184.2 ;
      RECT  184.6 202.0 192.2 202.8 ;
      RECT  191.4 200.4 192.2 202.0 ;
      RECT  189.6 196.8 190.4 197.2 ;
      RECT  186.2 192.8 187.8 193.6 ;
      RECT  189.6 198.0 190.4 200.4 ;
      RECT  184.6 194.2 192.2 195.0 ;
      RECT  189.4 201.2 190.2 202.0 ;
      RECT  188.4 195.0 189.2 195.2 ;
      RECT  187.2 200.4 188.2 201.2 ;
      RECT  184.6 195.6 185.4 199.8 ;
      RECT  187.2 199.8 188.0 200.4 ;
      RECT  184.6 200.4 185.4 202.0 ;
      RECT  189.2 197.2 190.4 198.0 ;
      RECT  189.0 192.8 190.6 193.6 ;
      RECT  189.6 196.0 190.6 196.8 ;
      RECT  189.4 200.4 190.4 201.2 ;
      RECT  187.0 196.0 188.0 196.8 ;
      RECT  187.2 196.8 188.0 199.0 ;
      RECT  187.2 199.0 188.8 199.8 ;
      RECT  191.4 195.6 192.2 199.8 ;
      RECT  184.6 202.8 192.2 202.0 ;
      RECT  191.4 204.4 192.2 202.8 ;
      RECT  189.6 208.0 190.4 207.6 ;
      RECT  186.2 212.0 187.8 211.2 ;
      RECT  189.6 206.8 190.4 204.4 ;
      RECT  184.6 210.6 192.2 209.8 ;
      RECT  189.4 203.6 190.2 202.8 ;
      RECT  188.4 209.8 189.2 209.6 ;
      RECT  187.2 204.4 188.2 203.6 ;
      RECT  184.6 209.2 185.4 205.0 ;
      RECT  187.2 205.0 188.0 204.4 ;
      RECT  184.6 204.4 185.4 202.8 ;
      RECT  189.2 207.6 190.4 206.8 ;
      RECT  189.0 212.0 190.6 211.2 ;
      RECT  189.6 208.8 190.6 208.0 ;
      RECT  189.4 204.4 190.4 203.6 ;
      RECT  187.0 208.8 188.0 208.0 ;
      RECT  187.2 208.0 188.0 205.8 ;
      RECT  187.2 205.8 188.8 205.0 ;
      RECT  191.4 209.2 192.2 205.0 ;
      RECT  184.6 222.8 192.2 223.6 ;
      RECT  191.4 221.2 192.2 222.8 ;
      RECT  189.6 217.6 190.4 218.0 ;
      RECT  186.2 213.6 187.8 214.4 ;
      RECT  189.6 218.8 190.4 221.2 ;
      RECT  184.6 215.0 192.2 215.8 ;
      RECT  189.4 222.0 190.2 222.8 ;
      RECT  188.4 215.8 189.2 216.0 ;
      RECT  187.2 221.2 188.2 222.0 ;
      RECT  184.6 216.4 185.4 220.6 ;
      RECT  187.2 220.6 188.0 221.2 ;
      RECT  184.6 221.2 185.4 222.8 ;
      RECT  189.2 218.0 190.4 218.8 ;
      RECT  189.0 213.6 190.6 214.4 ;
      RECT  189.6 216.8 190.6 217.6 ;
      RECT  189.4 221.2 190.4 222.0 ;
      RECT  187.0 216.8 188.0 217.6 ;
      RECT  187.2 217.6 188.0 219.8 ;
      RECT  187.2 219.8 188.8 220.6 ;
      RECT  191.4 216.4 192.2 220.6 ;
      RECT  184.6 223.6 192.2 222.8 ;
      RECT  191.4 225.2 192.2 223.6 ;
      RECT  189.6 228.8 190.4 228.4 ;
      RECT  186.2 232.8 187.8 232.0 ;
      RECT  189.6 227.6 190.4 225.2 ;
      RECT  184.6 231.4 192.2 230.6 ;
      RECT  189.4 224.4 190.2 223.6 ;
      RECT  188.4 230.6 189.2 230.4 ;
      RECT  187.2 225.2 188.2 224.4 ;
      RECT  184.6 230.0 185.4 225.8 ;
      RECT  187.2 225.8 188.0 225.2 ;
      RECT  184.6 225.2 185.4 223.6 ;
      RECT  189.2 228.4 190.4 227.6 ;
      RECT  189.0 232.8 190.6 232.0 ;
      RECT  189.6 229.6 190.6 228.8 ;
      RECT  189.4 225.2 190.4 224.4 ;
      RECT  187.0 229.6 188.0 228.8 ;
      RECT  187.2 228.8 188.0 226.6 ;
      RECT  187.2 226.6 188.8 225.8 ;
      RECT  191.4 230.0 192.2 225.8 ;
      RECT  184.6 243.6 192.2 244.4 ;
      RECT  191.4 242.0 192.2 243.6 ;
      RECT  189.6 238.4 190.4 238.8 ;
      RECT  186.2 234.4 187.8 235.2 ;
      RECT  189.6 239.6 190.4 242.0 ;
      RECT  184.6 235.8 192.2 236.6 ;
      RECT  189.4 242.8 190.2 243.6 ;
      RECT  188.4 236.6 189.2 236.8 ;
      RECT  187.2 242.0 188.2 242.8 ;
      RECT  184.6 237.2 185.4 241.4 ;
      RECT  187.2 241.4 188.0 242.0 ;
      RECT  184.6 242.0 185.4 243.6 ;
      RECT  189.2 238.8 190.4 239.6 ;
      RECT  189.0 234.4 190.6 235.2 ;
      RECT  189.6 237.6 190.6 238.4 ;
      RECT  189.4 242.0 190.4 242.8 ;
      RECT  187.0 237.6 188.0 238.4 ;
      RECT  187.2 238.4 188.0 240.6 ;
      RECT  187.2 240.6 188.8 241.4 ;
      RECT  191.4 237.2 192.2 241.4 ;
      RECT  184.6 244.4 192.2 243.6 ;
      RECT  191.4 246.0 192.2 244.4 ;
      RECT  189.6 249.6 190.4 249.2 ;
      RECT  186.2 253.6 187.8 252.8 ;
      RECT  189.6 248.4 190.4 246.0 ;
      RECT  184.6 252.2 192.2 251.4 ;
      RECT  189.4 245.2 190.2 244.4 ;
      RECT  188.4 251.4 189.2 251.2 ;
      RECT  187.2 246.0 188.2 245.2 ;
      RECT  184.6 250.8 185.4 246.6 ;
      RECT  187.2 246.6 188.0 246.0 ;
      RECT  184.6 246.0 185.4 244.4 ;
      RECT  189.2 249.2 190.4 248.4 ;
      RECT  189.0 253.6 190.6 252.8 ;
      RECT  189.6 250.4 190.6 249.6 ;
      RECT  189.4 246.0 190.4 245.2 ;
      RECT  187.0 250.4 188.0 249.6 ;
      RECT  187.2 249.6 188.0 247.4 ;
      RECT  187.2 247.4 188.8 246.6 ;
      RECT  191.4 250.8 192.2 246.6 ;
      RECT  184.6 264.4 192.2 265.2 ;
      RECT  191.4 262.8 192.2 264.4 ;
      RECT  189.6 259.2 190.4 259.6 ;
      RECT  186.2 255.2 187.8 256.0 ;
      RECT  189.6 260.4 190.4 262.8 ;
      RECT  184.6 256.6 192.2 257.4 ;
      RECT  189.4 263.6 190.2 264.4 ;
      RECT  188.4 257.4 189.2 257.6 ;
      RECT  187.2 262.8 188.2 263.6 ;
      RECT  184.6 258.0 185.4 262.2 ;
      RECT  187.2 262.2 188.0 262.8 ;
      RECT  184.6 262.8 185.4 264.4 ;
      RECT  189.2 259.6 190.4 260.4 ;
      RECT  189.0 255.2 190.6 256.0 ;
      RECT  189.6 258.4 190.6 259.2 ;
      RECT  189.4 262.8 190.4 263.6 ;
      RECT  187.0 258.4 188.0 259.2 ;
      RECT  187.2 259.2 188.0 261.4 ;
      RECT  187.2 261.4 188.8 262.2 ;
      RECT  191.4 258.0 192.2 262.2 ;
      RECT  184.6 265.2 192.2 264.4 ;
      RECT  191.4 266.8 192.2 265.2 ;
      RECT  189.6 270.4 190.4 270.0 ;
      RECT  186.2 274.4 187.8 273.6 ;
      RECT  189.6 269.2 190.4 266.8 ;
      RECT  184.6 273.0 192.2 272.2 ;
      RECT  189.4 266.0 190.2 265.2 ;
      RECT  188.4 272.2 189.2 272.0 ;
      RECT  187.2 266.8 188.2 266.0 ;
      RECT  184.6 271.6 185.4 267.4 ;
      RECT  187.2 267.4 188.0 266.8 ;
      RECT  184.6 266.8 185.4 265.2 ;
      RECT  189.2 270.0 190.4 269.2 ;
      RECT  189.0 274.4 190.6 273.6 ;
      RECT  189.6 271.2 190.6 270.4 ;
      RECT  189.4 266.8 190.4 266.0 ;
      RECT  187.0 271.2 188.0 270.4 ;
      RECT  187.2 270.4 188.0 268.2 ;
      RECT  187.2 268.2 188.8 267.4 ;
      RECT  191.4 271.6 192.2 267.4 ;
      RECT  184.6 285.2 192.2 286.0 ;
      RECT  191.4 283.6 192.2 285.2 ;
      RECT  189.6 280.0 190.4 280.4 ;
      RECT  186.2 276.0 187.8 276.8 ;
      RECT  189.6 281.2 190.4 283.6 ;
      RECT  184.6 277.4 192.2 278.2 ;
      RECT  189.4 284.4 190.2 285.2 ;
      RECT  188.4 278.2 189.2 278.4 ;
      RECT  187.2 283.6 188.2 284.4 ;
      RECT  184.6 278.8 185.4 283.0 ;
      RECT  187.2 283.0 188.0 283.6 ;
      RECT  184.6 283.6 185.4 285.2 ;
      RECT  189.2 280.4 190.4 281.2 ;
      RECT  189.0 276.0 190.6 276.8 ;
      RECT  189.6 279.2 190.6 280.0 ;
      RECT  189.4 283.6 190.4 284.4 ;
      RECT  187.0 279.2 188.0 280.0 ;
      RECT  187.2 280.0 188.0 282.2 ;
      RECT  187.2 282.2 188.8 283.0 ;
      RECT  191.4 278.8 192.2 283.0 ;
      RECT  184.6 286.0 192.2 285.2 ;
      RECT  191.4 287.6 192.2 286.0 ;
      RECT  189.6 291.2 190.4 290.8 ;
      RECT  186.2 295.2 187.8 294.4 ;
      RECT  189.6 290.0 190.4 287.6 ;
      RECT  184.6 293.8 192.2 293.0 ;
      RECT  189.4 286.8 190.2 286.0 ;
      RECT  188.4 293.0 189.2 292.8 ;
      RECT  187.2 287.6 188.2 286.8 ;
      RECT  184.6 292.4 185.4 288.2 ;
      RECT  187.2 288.2 188.0 287.6 ;
      RECT  184.6 287.6 185.4 286.0 ;
      RECT  189.2 290.8 190.4 290.0 ;
      RECT  189.0 295.2 190.6 294.4 ;
      RECT  189.6 292.0 190.6 291.2 ;
      RECT  189.4 287.6 190.4 286.8 ;
      RECT  187.0 292.0 188.0 291.2 ;
      RECT  187.2 291.2 188.0 289.0 ;
      RECT  187.2 289.0 188.8 288.2 ;
      RECT  191.4 292.4 192.2 288.2 ;
      RECT  184.6 306.0 192.2 306.8 ;
      RECT  191.4 304.4 192.2 306.0 ;
      RECT  189.6 300.8 190.4 301.2 ;
      RECT  186.2 296.8 187.8 297.6 ;
      RECT  189.6 302.0 190.4 304.4 ;
      RECT  184.6 298.2 192.2 299.0 ;
      RECT  189.4 305.2 190.2 306.0 ;
      RECT  188.4 299.0 189.2 299.2 ;
      RECT  187.2 304.4 188.2 305.2 ;
      RECT  184.6 299.6 185.4 303.8 ;
      RECT  187.2 303.8 188.0 304.4 ;
      RECT  184.6 304.4 185.4 306.0 ;
      RECT  189.2 301.2 190.4 302.0 ;
      RECT  189.0 296.8 190.6 297.6 ;
      RECT  189.6 300.0 190.6 300.8 ;
      RECT  189.4 304.4 190.4 305.2 ;
      RECT  187.0 300.0 188.0 300.8 ;
      RECT  187.2 300.8 188.0 303.0 ;
      RECT  187.2 303.0 188.8 303.8 ;
      RECT  191.4 299.6 192.2 303.8 ;
      RECT  184.6 306.8 192.2 306.0 ;
      RECT  191.4 308.4 192.2 306.8 ;
      RECT  189.6 312.0 190.4 311.6 ;
      RECT  186.2 316.0 187.8 315.2 ;
      RECT  189.6 310.8 190.4 308.4 ;
      RECT  184.6 314.6 192.2 313.8 ;
      RECT  189.4 307.6 190.2 306.8 ;
      RECT  188.4 313.8 189.2 313.6 ;
      RECT  187.2 308.4 188.2 307.6 ;
      RECT  184.6 313.2 185.4 309.0 ;
      RECT  187.2 309.0 188.0 308.4 ;
      RECT  184.6 308.4 185.4 306.8 ;
      RECT  189.2 311.6 190.4 310.8 ;
      RECT  189.0 316.0 190.6 315.2 ;
      RECT  189.6 312.8 190.6 312.0 ;
      RECT  189.4 308.4 190.4 307.6 ;
      RECT  187.0 312.8 188.0 312.0 ;
      RECT  187.2 312.0 188.0 309.8 ;
      RECT  187.2 309.8 188.8 309.0 ;
      RECT  191.4 313.2 192.2 309.0 ;
      RECT  184.6 326.8 192.2 327.6 ;
      RECT  191.4 325.2 192.2 326.8 ;
      RECT  189.6 321.6 190.4 322.0 ;
      RECT  186.2 317.6 187.8 318.4 ;
      RECT  189.6 322.8 190.4 325.2 ;
      RECT  184.6 319.0 192.2 319.8 ;
      RECT  189.4 326.0 190.2 326.8 ;
      RECT  188.4 319.8 189.2 320.0 ;
      RECT  187.2 325.2 188.2 326.0 ;
      RECT  184.6 320.4 185.4 324.6 ;
      RECT  187.2 324.6 188.0 325.2 ;
      RECT  184.6 325.2 185.4 326.8 ;
      RECT  189.2 322.0 190.4 322.8 ;
      RECT  189.0 317.6 190.6 318.4 ;
      RECT  189.6 320.8 190.6 321.6 ;
      RECT  189.4 325.2 190.4 326.0 ;
      RECT  187.0 320.8 188.0 321.6 ;
      RECT  187.2 321.6 188.0 323.8 ;
      RECT  187.2 323.8 188.8 324.6 ;
      RECT  191.4 320.4 192.2 324.6 ;
      RECT  184.6 327.6 192.2 326.8 ;
      RECT  191.4 329.2 192.2 327.6 ;
      RECT  189.6 332.8 190.4 332.4 ;
      RECT  186.2 336.8 187.8 336.0 ;
      RECT  189.6 331.6 190.4 329.2 ;
      RECT  184.6 335.4 192.2 334.6 ;
      RECT  189.4 328.4 190.2 327.6 ;
      RECT  188.4 334.6 189.2 334.4 ;
      RECT  187.2 329.2 188.2 328.4 ;
      RECT  184.6 334.0 185.4 329.8 ;
      RECT  187.2 329.8 188.0 329.2 ;
      RECT  184.6 329.2 185.4 327.6 ;
      RECT  189.2 332.4 190.4 331.6 ;
      RECT  189.0 336.8 190.6 336.0 ;
      RECT  189.6 333.6 190.6 332.8 ;
      RECT  189.4 329.2 190.4 328.4 ;
      RECT  187.0 333.6 188.0 332.8 ;
      RECT  187.2 332.8 188.0 330.6 ;
      RECT  187.2 330.6 188.8 329.8 ;
      RECT  191.4 334.0 192.2 329.8 ;
      RECT  184.6 347.6 192.2 348.4 ;
      RECT  191.4 346.0 192.2 347.6 ;
      RECT  189.6 342.4 190.4 342.8 ;
      RECT  186.2 338.4 187.8 339.2 ;
      RECT  189.6 343.6 190.4 346.0 ;
      RECT  184.6 339.8 192.2 340.6 ;
      RECT  189.4 346.8 190.2 347.6 ;
      RECT  188.4 340.6 189.2 340.8 ;
      RECT  187.2 346.0 188.2 346.8 ;
      RECT  184.6 341.2 185.4 345.4 ;
      RECT  187.2 345.4 188.0 346.0 ;
      RECT  184.6 346.0 185.4 347.6 ;
      RECT  189.2 342.8 190.4 343.6 ;
      RECT  189.0 338.4 190.6 339.2 ;
      RECT  189.6 341.6 190.6 342.4 ;
      RECT  189.4 346.0 190.4 346.8 ;
      RECT  187.0 341.6 188.0 342.4 ;
      RECT  187.2 342.4 188.0 344.6 ;
      RECT  187.2 344.6 188.8 345.4 ;
      RECT  191.4 341.2 192.2 345.4 ;
      RECT  184.6 348.4 192.2 347.6 ;
      RECT  191.4 350.0 192.2 348.4 ;
      RECT  189.6 353.6 190.4 353.2 ;
      RECT  186.2 357.6 187.8 356.8 ;
      RECT  189.6 352.4 190.4 350.0 ;
      RECT  184.6 356.2 192.2 355.4 ;
      RECT  189.4 349.2 190.2 348.4 ;
      RECT  188.4 355.4 189.2 355.2 ;
      RECT  187.2 350.0 188.2 349.2 ;
      RECT  184.6 354.8 185.4 350.6 ;
      RECT  187.2 350.6 188.0 350.0 ;
      RECT  184.6 350.0 185.4 348.4 ;
      RECT  189.2 353.2 190.4 352.4 ;
      RECT  189.0 357.6 190.6 356.8 ;
      RECT  189.6 354.4 190.6 353.6 ;
      RECT  189.4 350.0 190.4 349.2 ;
      RECT  187.0 354.4 188.0 353.6 ;
      RECT  187.2 353.6 188.0 351.4 ;
      RECT  187.2 351.4 188.8 350.6 ;
      RECT  191.4 354.8 192.2 350.6 ;
      RECT  184.6 368.4 192.2 369.2 ;
      RECT  191.4 366.8 192.2 368.4 ;
      RECT  189.6 363.2 190.4 363.6 ;
      RECT  189.6 364.4 190.4 366.8 ;
      RECT  184.6 360.6 192.2 361.4 ;
      RECT  189.8 359.2 190.6 360.0 ;
      RECT  188.4 361.4 189.2 361.6 ;
      RECT  187.2 366.8 188.2 367.6 ;
      RECT  184.6 362.0 185.4 366.2 ;
      RECT  187.2 366.2 188.0 366.8 ;
      RECT  184.6 366.8 185.4 368.4 ;
      RECT  189.2 363.6 190.4 364.4 ;
      RECT  189.6 362.4 190.6 363.2 ;
      RECT  189.4 366.8 190.4 367.6 ;
      RECT  187.0 362.4 188.0 363.2 ;
      RECT  187.2 363.2 188.0 365.4 ;
      RECT  187.2 365.4 188.8 366.2 ;
      RECT  187.0 359.2 187.8 360.0 ;
      RECT  191.4 362.0 192.2 366.2 ;
      RECT  185.0 173.4 191.8 174.2 ;
      RECT  185.0 189.0 191.8 189.8 ;
      RECT  185.0 194.2 191.8 195.0 ;
      RECT  185.0 209.8 191.8 210.6 ;
      RECT  185.0 215.0 191.8 215.8 ;
      RECT  185.0 230.6 191.8 231.4 ;
      RECT  185.0 235.8 191.8 236.6 ;
      RECT  185.0 251.4 191.8 252.2 ;
      RECT  185.0 256.6 191.8 257.4 ;
      RECT  185.0 272.2 191.8 273.0 ;
      RECT  185.0 277.4 191.8 278.2 ;
      RECT  185.0 293.0 191.8 293.8 ;
      RECT  185.0 298.2 191.8 299.0 ;
      RECT  185.0 313.8 191.8 314.6 ;
      RECT  185.0 319.0 191.8 319.8 ;
      RECT  185.0 334.6 191.8 335.4 ;
      RECT  185.0 339.8 191.8 340.6 ;
      RECT  185.0 355.4 191.8 356.2 ;
      RECT  185.0 360.6 191.8 361.4 ;
      RECT  191.4 182.0 199.0 181.2 ;
      RECT  198.2 183.6 199.0 182.0 ;
      RECT  196.4 187.2 197.2 186.8 ;
      RECT  196.4 186.0 197.2 183.6 ;
      RECT  191.4 189.8 199.0 189.0 ;
      RECT  196.6 191.2 197.4 190.4 ;
      RECT  195.2 189.0 196.0 188.8 ;
      RECT  194.0 183.6 195.0 182.8 ;
      RECT  191.4 188.4 192.2 184.2 ;
      RECT  194.0 184.2 194.8 183.6 ;
      RECT  191.4 183.6 192.2 182.0 ;
      RECT  196.0 186.8 197.2 186.0 ;
      RECT  196.4 188.0 197.4 187.2 ;
      RECT  196.2 183.6 197.2 182.8 ;
      RECT  193.8 188.0 194.8 187.2 ;
      RECT  194.0 187.2 194.8 185.0 ;
      RECT  194.0 185.0 195.6 184.2 ;
      RECT  193.8 191.2 194.6 190.4 ;
      RECT  198.2 188.4 199.0 184.2 ;
      RECT  198.2 182.0 205.8 181.2 ;
      RECT  205.0 183.6 205.8 182.0 ;
      RECT  203.2 187.2 204.0 186.8 ;
      RECT  203.2 186.0 204.0 183.6 ;
      RECT  198.2 189.8 205.8 189.0 ;
      RECT  203.4 191.2 204.2 190.4 ;
      RECT  202.0 189.0 202.8 188.8 ;
      RECT  200.8 183.6 201.8 182.8 ;
      RECT  198.2 188.4 199.0 184.2 ;
      RECT  200.8 184.2 201.6 183.6 ;
      RECT  198.2 183.6 199.0 182.0 ;
      RECT  202.8 186.8 204.0 186.0 ;
      RECT  203.2 188.0 204.2 187.2 ;
      RECT  203.0 183.6 204.0 182.8 ;
      RECT  200.6 188.0 201.6 187.2 ;
      RECT  200.8 187.2 201.6 185.0 ;
      RECT  200.8 185.0 202.4 184.2 ;
      RECT  200.6 191.2 201.4 190.4 ;
      RECT  205.0 188.4 205.8 184.2 ;
      RECT  191.8 189.8 205.4 189.0 ;
      RECT  191.4 181.2 199.0 182.0 ;
      RECT  198.2 179.6 199.0 181.2 ;
      RECT  196.4 176.0 197.2 176.4 ;
      RECT  196.4 177.2 197.2 179.6 ;
      RECT  191.4 173.4 199.0 174.2 ;
      RECT  196.6 172.0 197.4 172.8 ;
      RECT  195.2 174.2 196.0 174.4 ;
      RECT  194.0 179.6 195.0 180.4 ;
      RECT  191.4 174.8 192.2 179.0 ;
      RECT  194.0 179.0 194.8 179.6 ;
      RECT  191.4 179.6 192.2 181.2 ;
      RECT  196.0 176.4 197.2 177.2 ;
      RECT  196.4 175.2 197.4 176.0 ;
      RECT  196.2 179.6 197.2 180.4 ;
      RECT  193.8 175.2 194.8 176.0 ;
      RECT  194.0 176.0 194.8 178.2 ;
      RECT  194.0 178.2 195.6 179.0 ;
      RECT  193.8 172.0 194.6 172.8 ;
      RECT  198.2 174.8 199.0 179.0 ;
      RECT  198.2 181.2 205.8 182.0 ;
      RECT  205.0 179.6 205.8 181.2 ;
      RECT  203.2 176.0 204.0 176.4 ;
      RECT  203.2 177.2 204.0 179.6 ;
      RECT  198.2 173.4 205.8 174.2 ;
      RECT  203.4 172.0 204.2 172.8 ;
      RECT  202.0 174.2 202.8 174.4 ;
      RECT  200.8 179.6 201.8 180.4 ;
      RECT  198.2 174.8 199.0 179.0 ;
      RECT  200.8 179.0 201.6 179.6 ;
      RECT  198.2 179.6 199.0 181.2 ;
      RECT  202.8 176.4 204.0 177.2 ;
      RECT  203.2 175.2 204.2 176.0 ;
      RECT  203.0 179.6 204.0 180.4 ;
      RECT  200.6 175.2 201.6 176.0 ;
      RECT  200.8 176.0 201.6 178.2 ;
      RECT  200.8 178.2 202.4 179.0 ;
      RECT  200.6 172.0 201.4 172.8 ;
      RECT  205.0 174.8 205.8 179.0 ;
      RECT  191.8 173.4 205.4 174.2 ;
      RECT  191.4 368.4 199.0 369.2 ;
      RECT  198.2 366.8 199.0 368.4 ;
      RECT  196.4 363.2 197.2 363.6 ;
      RECT  196.4 364.4 197.2 366.8 ;
      RECT  191.4 360.6 199.0 361.4 ;
      RECT  196.6 359.2 197.4 360.0 ;
      RECT  195.2 361.4 196.0 361.6 ;
      RECT  194.0 366.8 195.0 367.6 ;
      RECT  191.4 362.0 192.2 366.2 ;
      RECT  194.0 366.2 194.8 366.8 ;
      RECT  191.4 366.8 192.2 368.4 ;
      RECT  196.0 363.6 197.2 364.4 ;
      RECT  196.4 362.4 197.4 363.2 ;
      RECT  196.2 366.8 197.2 367.6 ;
      RECT  193.8 362.4 194.8 363.2 ;
      RECT  194.0 363.2 194.8 365.4 ;
      RECT  194.0 365.4 195.6 366.2 ;
      RECT  193.8 359.2 194.6 360.0 ;
      RECT  198.2 362.0 199.0 366.2 ;
      RECT  198.2 368.4 205.8 369.2 ;
      RECT  205.0 366.8 205.8 368.4 ;
      RECT  203.2 363.2 204.0 363.6 ;
      RECT  203.2 364.4 204.0 366.8 ;
      RECT  198.2 360.6 205.8 361.4 ;
      RECT  203.4 359.2 204.2 360.0 ;
      RECT  202.0 361.4 202.8 361.6 ;
      RECT  200.8 366.8 201.8 367.6 ;
      RECT  198.2 362.0 199.0 366.2 ;
      RECT  200.8 366.2 201.6 366.8 ;
      RECT  198.2 366.8 199.0 368.4 ;
      RECT  202.8 363.6 204.0 364.4 ;
      RECT  203.2 362.4 204.2 363.2 ;
      RECT  203.0 366.8 204.0 367.6 ;
      RECT  200.6 362.4 201.6 363.2 ;
      RECT  200.8 363.2 201.6 365.4 ;
      RECT  200.8 365.4 202.4 366.2 ;
      RECT  200.6 359.2 201.4 360.0 ;
      RECT  205.0 362.0 205.8 366.2 ;
      RECT  191.8 360.6 205.4 361.4 ;
      RECT  177.8 181.2 185.4 182.0 ;
      RECT  184.6 179.6 185.4 181.2 ;
      RECT  182.8 176.0 183.6 176.4 ;
      RECT  182.8 177.2 183.6 179.6 ;
      RECT  177.8 173.4 185.4 174.2 ;
      RECT  183.0 172.0 183.8 172.8 ;
      RECT  181.6 174.2 182.4 174.4 ;
      RECT  180.4 179.6 181.4 180.4 ;
      RECT  177.8 174.8 178.6 179.0 ;
      RECT  180.4 179.0 181.2 179.6 ;
      RECT  177.8 179.6 178.6 181.2 ;
      RECT  182.4 176.4 183.6 177.2 ;
      RECT  182.8 175.2 183.8 176.0 ;
      RECT  182.6 179.6 183.6 180.4 ;
      RECT  180.2 175.2 181.2 176.0 ;
      RECT  180.4 176.0 181.2 178.2 ;
      RECT  180.4 178.2 182.0 179.0 ;
      RECT  180.2 172.0 181.0 172.8 ;
      RECT  184.6 174.8 185.4 179.0 ;
      RECT  177.8 182.0 185.4 181.2 ;
      RECT  184.6 183.6 185.4 182.0 ;
      RECT  182.8 187.2 183.6 186.8 ;
      RECT  182.8 186.0 183.6 183.6 ;
      RECT  177.8 189.8 185.4 189.0 ;
      RECT  183.0 191.2 183.8 190.4 ;
      RECT  181.6 189.0 182.4 188.8 ;
      RECT  180.4 183.6 181.4 182.8 ;
      RECT  177.8 188.4 178.6 184.2 ;
      RECT  180.4 184.2 181.2 183.6 ;
      RECT  177.8 183.6 178.6 182.0 ;
      RECT  182.4 186.8 183.6 186.0 ;
      RECT  182.8 188.0 183.8 187.2 ;
      RECT  182.6 183.6 183.6 182.8 ;
      RECT  180.2 188.0 181.2 187.2 ;
      RECT  180.4 187.2 181.2 185.0 ;
      RECT  180.4 185.0 182.0 184.2 ;
      RECT  180.2 191.2 181.0 190.4 ;
      RECT  184.6 188.4 185.4 184.2 ;
      RECT  177.8 202.0 185.4 202.8 ;
      RECT  184.6 200.4 185.4 202.0 ;
      RECT  182.8 196.8 183.6 197.2 ;
      RECT  182.8 198.0 183.6 200.4 ;
      RECT  177.8 194.2 185.4 195.0 ;
      RECT  183.0 192.8 183.8 193.6 ;
      RECT  181.6 195.0 182.4 195.2 ;
      RECT  180.4 200.4 181.4 201.2 ;
      RECT  177.8 195.6 178.6 199.8 ;
      RECT  180.4 199.8 181.2 200.4 ;
      RECT  177.8 200.4 178.6 202.0 ;
      RECT  182.4 197.2 183.6 198.0 ;
      RECT  182.8 196.0 183.8 196.8 ;
      RECT  182.6 200.4 183.6 201.2 ;
      RECT  180.2 196.0 181.2 196.8 ;
      RECT  180.4 196.8 181.2 199.0 ;
      RECT  180.4 199.0 182.0 199.8 ;
      RECT  180.2 192.8 181.0 193.6 ;
      RECT  184.6 195.6 185.4 199.8 ;
      RECT  177.8 202.8 185.4 202.0 ;
      RECT  184.6 204.4 185.4 202.8 ;
      RECT  182.8 208.0 183.6 207.6 ;
      RECT  182.8 206.8 183.6 204.4 ;
      RECT  177.8 210.6 185.4 209.8 ;
      RECT  183.0 212.0 183.8 211.2 ;
      RECT  181.6 209.8 182.4 209.6 ;
      RECT  180.4 204.4 181.4 203.6 ;
      RECT  177.8 209.2 178.6 205.0 ;
      RECT  180.4 205.0 181.2 204.4 ;
      RECT  177.8 204.4 178.6 202.8 ;
      RECT  182.4 207.6 183.6 206.8 ;
      RECT  182.8 208.8 183.8 208.0 ;
      RECT  182.6 204.4 183.6 203.6 ;
      RECT  180.2 208.8 181.2 208.0 ;
      RECT  180.4 208.0 181.2 205.8 ;
      RECT  180.4 205.8 182.0 205.0 ;
      RECT  180.2 212.0 181.0 211.2 ;
      RECT  184.6 209.2 185.4 205.0 ;
      RECT  177.8 222.8 185.4 223.6 ;
      RECT  184.6 221.2 185.4 222.8 ;
      RECT  182.8 217.6 183.6 218.0 ;
      RECT  182.8 218.8 183.6 221.2 ;
      RECT  177.8 215.0 185.4 215.8 ;
      RECT  183.0 213.6 183.8 214.4 ;
      RECT  181.6 215.8 182.4 216.0 ;
      RECT  180.4 221.2 181.4 222.0 ;
      RECT  177.8 216.4 178.6 220.6 ;
      RECT  180.4 220.6 181.2 221.2 ;
      RECT  177.8 221.2 178.6 222.8 ;
      RECT  182.4 218.0 183.6 218.8 ;
      RECT  182.8 216.8 183.8 217.6 ;
      RECT  182.6 221.2 183.6 222.0 ;
      RECT  180.2 216.8 181.2 217.6 ;
      RECT  180.4 217.6 181.2 219.8 ;
      RECT  180.4 219.8 182.0 220.6 ;
      RECT  180.2 213.6 181.0 214.4 ;
      RECT  184.6 216.4 185.4 220.6 ;
      RECT  177.8 223.6 185.4 222.8 ;
      RECT  184.6 225.2 185.4 223.6 ;
      RECT  182.8 228.8 183.6 228.4 ;
      RECT  182.8 227.6 183.6 225.2 ;
      RECT  177.8 231.4 185.4 230.6 ;
      RECT  183.0 232.8 183.8 232.0 ;
      RECT  181.6 230.6 182.4 230.4 ;
      RECT  180.4 225.2 181.4 224.4 ;
      RECT  177.8 230.0 178.6 225.8 ;
      RECT  180.4 225.8 181.2 225.2 ;
      RECT  177.8 225.2 178.6 223.6 ;
      RECT  182.4 228.4 183.6 227.6 ;
      RECT  182.8 229.6 183.8 228.8 ;
      RECT  182.6 225.2 183.6 224.4 ;
      RECT  180.2 229.6 181.2 228.8 ;
      RECT  180.4 228.8 181.2 226.6 ;
      RECT  180.4 226.6 182.0 225.8 ;
      RECT  180.2 232.8 181.0 232.0 ;
      RECT  184.6 230.0 185.4 225.8 ;
      RECT  177.8 243.6 185.4 244.4 ;
      RECT  184.6 242.0 185.4 243.6 ;
      RECT  182.8 238.4 183.6 238.8 ;
      RECT  182.8 239.6 183.6 242.0 ;
      RECT  177.8 235.8 185.4 236.6 ;
      RECT  183.0 234.4 183.8 235.2 ;
      RECT  181.6 236.6 182.4 236.8 ;
      RECT  180.4 242.0 181.4 242.8 ;
      RECT  177.8 237.2 178.6 241.4 ;
      RECT  180.4 241.4 181.2 242.0 ;
      RECT  177.8 242.0 178.6 243.6 ;
      RECT  182.4 238.8 183.6 239.6 ;
      RECT  182.8 237.6 183.8 238.4 ;
      RECT  182.6 242.0 183.6 242.8 ;
      RECT  180.2 237.6 181.2 238.4 ;
      RECT  180.4 238.4 181.2 240.6 ;
      RECT  180.4 240.6 182.0 241.4 ;
      RECT  180.2 234.4 181.0 235.2 ;
      RECT  184.6 237.2 185.4 241.4 ;
      RECT  177.8 244.4 185.4 243.6 ;
      RECT  184.6 246.0 185.4 244.4 ;
      RECT  182.8 249.6 183.6 249.2 ;
      RECT  182.8 248.4 183.6 246.0 ;
      RECT  177.8 252.2 185.4 251.4 ;
      RECT  183.0 253.6 183.8 252.8 ;
      RECT  181.6 251.4 182.4 251.2 ;
      RECT  180.4 246.0 181.4 245.2 ;
      RECT  177.8 250.8 178.6 246.6 ;
      RECT  180.4 246.6 181.2 246.0 ;
      RECT  177.8 246.0 178.6 244.4 ;
      RECT  182.4 249.2 183.6 248.4 ;
      RECT  182.8 250.4 183.8 249.6 ;
      RECT  182.6 246.0 183.6 245.2 ;
      RECT  180.2 250.4 181.2 249.6 ;
      RECT  180.4 249.6 181.2 247.4 ;
      RECT  180.4 247.4 182.0 246.6 ;
      RECT  180.2 253.6 181.0 252.8 ;
      RECT  184.6 250.8 185.4 246.6 ;
      RECT  177.8 264.4 185.4 265.2 ;
      RECT  184.6 262.8 185.4 264.4 ;
      RECT  182.8 259.2 183.6 259.6 ;
      RECT  182.8 260.4 183.6 262.8 ;
      RECT  177.8 256.6 185.4 257.4 ;
      RECT  183.0 255.2 183.8 256.0 ;
      RECT  181.6 257.4 182.4 257.6 ;
      RECT  180.4 262.8 181.4 263.6 ;
      RECT  177.8 258.0 178.6 262.2 ;
      RECT  180.4 262.2 181.2 262.8 ;
      RECT  177.8 262.8 178.6 264.4 ;
      RECT  182.4 259.6 183.6 260.4 ;
      RECT  182.8 258.4 183.8 259.2 ;
      RECT  182.6 262.8 183.6 263.6 ;
      RECT  180.2 258.4 181.2 259.2 ;
      RECT  180.4 259.2 181.2 261.4 ;
      RECT  180.4 261.4 182.0 262.2 ;
      RECT  180.2 255.2 181.0 256.0 ;
      RECT  184.6 258.0 185.4 262.2 ;
      RECT  177.8 265.2 185.4 264.4 ;
      RECT  184.6 266.8 185.4 265.2 ;
      RECT  182.8 270.4 183.6 270.0 ;
      RECT  182.8 269.2 183.6 266.8 ;
      RECT  177.8 273.0 185.4 272.2 ;
      RECT  183.0 274.4 183.8 273.6 ;
      RECT  181.6 272.2 182.4 272.0 ;
      RECT  180.4 266.8 181.4 266.0 ;
      RECT  177.8 271.6 178.6 267.4 ;
      RECT  180.4 267.4 181.2 266.8 ;
      RECT  177.8 266.8 178.6 265.2 ;
      RECT  182.4 270.0 183.6 269.2 ;
      RECT  182.8 271.2 183.8 270.4 ;
      RECT  182.6 266.8 183.6 266.0 ;
      RECT  180.2 271.2 181.2 270.4 ;
      RECT  180.4 270.4 181.2 268.2 ;
      RECT  180.4 268.2 182.0 267.4 ;
      RECT  180.2 274.4 181.0 273.6 ;
      RECT  184.6 271.6 185.4 267.4 ;
      RECT  177.8 285.2 185.4 286.0 ;
      RECT  184.6 283.6 185.4 285.2 ;
      RECT  182.8 280.0 183.6 280.4 ;
      RECT  182.8 281.2 183.6 283.6 ;
      RECT  177.8 277.4 185.4 278.2 ;
      RECT  183.0 276.0 183.8 276.8 ;
      RECT  181.6 278.2 182.4 278.4 ;
      RECT  180.4 283.6 181.4 284.4 ;
      RECT  177.8 278.8 178.6 283.0 ;
      RECT  180.4 283.0 181.2 283.6 ;
      RECT  177.8 283.6 178.6 285.2 ;
      RECT  182.4 280.4 183.6 281.2 ;
      RECT  182.8 279.2 183.8 280.0 ;
      RECT  182.6 283.6 183.6 284.4 ;
      RECT  180.2 279.2 181.2 280.0 ;
      RECT  180.4 280.0 181.2 282.2 ;
      RECT  180.4 282.2 182.0 283.0 ;
      RECT  180.2 276.0 181.0 276.8 ;
      RECT  184.6 278.8 185.4 283.0 ;
      RECT  177.8 286.0 185.4 285.2 ;
      RECT  184.6 287.6 185.4 286.0 ;
      RECT  182.8 291.2 183.6 290.8 ;
      RECT  182.8 290.0 183.6 287.6 ;
      RECT  177.8 293.8 185.4 293.0 ;
      RECT  183.0 295.2 183.8 294.4 ;
      RECT  181.6 293.0 182.4 292.8 ;
      RECT  180.4 287.6 181.4 286.8 ;
      RECT  177.8 292.4 178.6 288.2 ;
      RECT  180.4 288.2 181.2 287.6 ;
      RECT  177.8 287.6 178.6 286.0 ;
      RECT  182.4 290.8 183.6 290.0 ;
      RECT  182.8 292.0 183.8 291.2 ;
      RECT  182.6 287.6 183.6 286.8 ;
      RECT  180.2 292.0 181.2 291.2 ;
      RECT  180.4 291.2 181.2 289.0 ;
      RECT  180.4 289.0 182.0 288.2 ;
      RECT  180.2 295.2 181.0 294.4 ;
      RECT  184.6 292.4 185.4 288.2 ;
      RECT  177.8 306.0 185.4 306.8 ;
      RECT  184.6 304.4 185.4 306.0 ;
      RECT  182.8 300.8 183.6 301.2 ;
      RECT  182.8 302.0 183.6 304.4 ;
      RECT  177.8 298.2 185.4 299.0 ;
      RECT  183.0 296.8 183.8 297.6 ;
      RECT  181.6 299.0 182.4 299.2 ;
      RECT  180.4 304.4 181.4 305.2 ;
      RECT  177.8 299.6 178.6 303.8 ;
      RECT  180.4 303.8 181.2 304.4 ;
      RECT  177.8 304.4 178.6 306.0 ;
      RECT  182.4 301.2 183.6 302.0 ;
      RECT  182.8 300.0 183.8 300.8 ;
      RECT  182.6 304.4 183.6 305.2 ;
      RECT  180.2 300.0 181.2 300.8 ;
      RECT  180.4 300.8 181.2 303.0 ;
      RECT  180.4 303.0 182.0 303.8 ;
      RECT  180.2 296.8 181.0 297.6 ;
      RECT  184.6 299.6 185.4 303.8 ;
      RECT  177.8 306.8 185.4 306.0 ;
      RECT  184.6 308.4 185.4 306.8 ;
      RECT  182.8 312.0 183.6 311.6 ;
      RECT  182.8 310.8 183.6 308.4 ;
      RECT  177.8 314.6 185.4 313.8 ;
      RECT  183.0 316.0 183.8 315.2 ;
      RECT  181.6 313.8 182.4 313.6 ;
      RECT  180.4 308.4 181.4 307.6 ;
      RECT  177.8 313.2 178.6 309.0 ;
      RECT  180.4 309.0 181.2 308.4 ;
      RECT  177.8 308.4 178.6 306.8 ;
      RECT  182.4 311.6 183.6 310.8 ;
      RECT  182.8 312.8 183.8 312.0 ;
      RECT  182.6 308.4 183.6 307.6 ;
      RECT  180.2 312.8 181.2 312.0 ;
      RECT  180.4 312.0 181.2 309.8 ;
      RECT  180.4 309.8 182.0 309.0 ;
      RECT  180.2 316.0 181.0 315.2 ;
      RECT  184.6 313.2 185.4 309.0 ;
      RECT  177.8 326.8 185.4 327.6 ;
      RECT  184.6 325.2 185.4 326.8 ;
      RECT  182.8 321.6 183.6 322.0 ;
      RECT  182.8 322.8 183.6 325.2 ;
      RECT  177.8 319.0 185.4 319.8 ;
      RECT  183.0 317.6 183.8 318.4 ;
      RECT  181.6 319.8 182.4 320.0 ;
      RECT  180.4 325.2 181.4 326.0 ;
      RECT  177.8 320.4 178.6 324.6 ;
      RECT  180.4 324.6 181.2 325.2 ;
      RECT  177.8 325.2 178.6 326.8 ;
      RECT  182.4 322.0 183.6 322.8 ;
      RECT  182.8 320.8 183.8 321.6 ;
      RECT  182.6 325.2 183.6 326.0 ;
      RECT  180.2 320.8 181.2 321.6 ;
      RECT  180.4 321.6 181.2 323.8 ;
      RECT  180.4 323.8 182.0 324.6 ;
      RECT  180.2 317.6 181.0 318.4 ;
      RECT  184.6 320.4 185.4 324.6 ;
      RECT  177.8 327.6 185.4 326.8 ;
      RECT  184.6 329.2 185.4 327.6 ;
      RECT  182.8 332.8 183.6 332.4 ;
      RECT  182.8 331.6 183.6 329.2 ;
      RECT  177.8 335.4 185.4 334.6 ;
      RECT  183.0 336.8 183.8 336.0 ;
      RECT  181.6 334.6 182.4 334.4 ;
      RECT  180.4 329.2 181.4 328.4 ;
      RECT  177.8 334.0 178.6 329.8 ;
      RECT  180.4 329.8 181.2 329.2 ;
      RECT  177.8 329.2 178.6 327.6 ;
      RECT  182.4 332.4 183.6 331.6 ;
      RECT  182.8 333.6 183.8 332.8 ;
      RECT  182.6 329.2 183.6 328.4 ;
      RECT  180.2 333.6 181.2 332.8 ;
      RECT  180.4 332.8 181.2 330.6 ;
      RECT  180.4 330.6 182.0 329.8 ;
      RECT  180.2 336.8 181.0 336.0 ;
      RECT  184.6 334.0 185.4 329.8 ;
      RECT  177.8 347.6 185.4 348.4 ;
      RECT  184.6 346.0 185.4 347.6 ;
      RECT  182.8 342.4 183.6 342.8 ;
      RECT  182.8 343.6 183.6 346.0 ;
      RECT  177.8 339.8 185.4 340.6 ;
      RECT  183.0 338.4 183.8 339.2 ;
      RECT  181.6 340.6 182.4 340.8 ;
      RECT  180.4 346.0 181.4 346.8 ;
      RECT  177.8 341.2 178.6 345.4 ;
      RECT  180.4 345.4 181.2 346.0 ;
      RECT  177.8 346.0 178.6 347.6 ;
      RECT  182.4 342.8 183.6 343.6 ;
      RECT  182.8 341.6 183.8 342.4 ;
      RECT  182.6 346.0 183.6 346.8 ;
      RECT  180.2 341.6 181.2 342.4 ;
      RECT  180.4 342.4 181.2 344.6 ;
      RECT  180.4 344.6 182.0 345.4 ;
      RECT  180.2 338.4 181.0 339.2 ;
      RECT  184.6 341.2 185.4 345.4 ;
      RECT  177.8 348.4 185.4 347.6 ;
      RECT  184.6 350.0 185.4 348.4 ;
      RECT  182.8 353.6 183.6 353.2 ;
      RECT  182.8 352.4 183.6 350.0 ;
      RECT  177.8 356.2 185.4 355.4 ;
      RECT  183.0 357.6 183.8 356.8 ;
      RECT  181.6 355.4 182.4 355.2 ;
      RECT  180.4 350.0 181.4 349.2 ;
      RECT  177.8 354.8 178.6 350.6 ;
      RECT  180.4 350.6 181.2 350.0 ;
      RECT  177.8 350.0 178.6 348.4 ;
      RECT  182.4 353.2 183.6 352.4 ;
      RECT  182.8 354.4 183.8 353.6 ;
      RECT  182.6 350.0 183.6 349.2 ;
      RECT  180.2 354.4 181.2 353.6 ;
      RECT  180.4 353.6 181.2 351.4 ;
      RECT  180.4 351.4 182.0 350.6 ;
      RECT  180.2 357.6 181.0 356.8 ;
      RECT  184.6 354.8 185.4 350.6 ;
      RECT  177.8 368.4 185.4 369.2 ;
      RECT  184.6 366.8 185.4 368.4 ;
      RECT  182.8 363.2 183.6 363.6 ;
      RECT  182.8 364.4 183.6 366.8 ;
      RECT  177.8 360.6 185.4 361.4 ;
      RECT  183.0 359.2 183.8 360.0 ;
      RECT  181.6 361.4 182.4 361.6 ;
      RECT  180.4 366.8 181.4 367.6 ;
      RECT  177.8 362.0 178.6 366.2 ;
      RECT  180.4 366.2 181.2 366.8 ;
      RECT  177.8 366.8 178.6 368.4 ;
      RECT  182.4 363.6 183.6 364.4 ;
      RECT  182.8 362.4 183.8 363.2 ;
      RECT  182.6 366.8 183.6 367.6 ;
      RECT  180.2 362.4 181.2 363.2 ;
      RECT  180.4 363.2 181.2 365.4 ;
      RECT  180.4 365.4 182.0 366.2 ;
      RECT  180.2 359.2 181.0 360.0 ;
      RECT  184.6 362.0 185.4 366.2 ;
      RECT  178.2 173.4 185.0 174.2 ;
      RECT  178.2 189.0 185.0 189.8 ;
      RECT  178.2 194.2 185.0 195.0 ;
      RECT  178.2 209.8 185.0 210.6 ;
      RECT  178.2 215.0 185.0 215.8 ;
      RECT  178.2 230.6 185.0 231.4 ;
      RECT  178.2 235.8 185.0 236.6 ;
      RECT  178.2 251.4 185.0 252.2 ;
      RECT  178.2 256.6 185.0 257.4 ;
      RECT  178.2 272.2 185.0 273.0 ;
      RECT  178.2 277.4 185.0 278.2 ;
      RECT  178.2 293.0 185.0 293.8 ;
      RECT  178.2 298.2 185.0 299.0 ;
      RECT  178.2 313.8 185.0 314.6 ;
      RECT  178.2 319.0 185.0 319.8 ;
      RECT  178.2 334.6 185.0 335.4 ;
      RECT  178.2 339.8 185.0 340.6 ;
      RECT  178.2 355.4 185.0 356.2 ;
      RECT  178.2 360.6 185.0 361.4 ;
      RECT  205.0 181.2 212.6 182.0 ;
      RECT  211.8 179.6 212.6 181.2 ;
      RECT  210.0 176.0 210.8 176.4 ;
      RECT  210.0 177.2 210.8 179.6 ;
      RECT  205.0 173.4 212.6 174.2 ;
      RECT  210.2 172.0 211.0 172.8 ;
      RECT  208.8 174.2 209.6 174.4 ;
      RECT  207.6 179.6 208.6 180.4 ;
      RECT  205.0 174.8 205.8 179.0 ;
      RECT  207.6 179.0 208.4 179.6 ;
      RECT  205.0 179.6 205.8 181.2 ;
      RECT  209.6 176.4 210.8 177.2 ;
      RECT  210.0 175.2 211.0 176.0 ;
      RECT  209.8 179.6 210.8 180.4 ;
      RECT  207.4 175.2 208.4 176.0 ;
      RECT  207.6 176.0 208.4 178.2 ;
      RECT  207.6 178.2 209.2 179.0 ;
      RECT  207.4 172.0 208.2 172.8 ;
      RECT  211.8 174.8 212.6 179.0 ;
      RECT  205.0 182.0 212.6 181.2 ;
      RECT  211.8 183.6 212.6 182.0 ;
      RECT  210.0 187.2 210.8 186.8 ;
      RECT  210.0 186.0 210.8 183.6 ;
      RECT  205.0 189.8 212.6 189.0 ;
      RECT  210.2 191.2 211.0 190.4 ;
      RECT  208.8 189.0 209.6 188.8 ;
      RECT  207.6 183.6 208.6 182.8 ;
      RECT  205.0 188.4 205.8 184.2 ;
      RECT  207.6 184.2 208.4 183.6 ;
      RECT  205.0 183.6 205.8 182.0 ;
      RECT  209.6 186.8 210.8 186.0 ;
      RECT  210.0 188.0 211.0 187.2 ;
      RECT  209.8 183.6 210.8 182.8 ;
      RECT  207.4 188.0 208.4 187.2 ;
      RECT  207.6 187.2 208.4 185.0 ;
      RECT  207.6 185.0 209.2 184.2 ;
      RECT  207.4 191.2 208.2 190.4 ;
      RECT  211.8 188.4 212.6 184.2 ;
      RECT  205.0 202.0 212.6 202.8 ;
      RECT  211.8 200.4 212.6 202.0 ;
      RECT  210.0 196.8 210.8 197.2 ;
      RECT  210.0 198.0 210.8 200.4 ;
      RECT  205.0 194.2 212.6 195.0 ;
      RECT  210.2 192.8 211.0 193.6 ;
      RECT  208.8 195.0 209.6 195.2 ;
      RECT  207.6 200.4 208.6 201.2 ;
      RECT  205.0 195.6 205.8 199.8 ;
      RECT  207.6 199.8 208.4 200.4 ;
      RECT  205.0 200.4 205.8 202.0 ;
      RECT  209.6 197.2 210.8 198.0 ;
      RECT  210.0 196.0 211.0 196.8 ;
      RECT  209.8 200.4 210.8 201.2 ;
      RECT  207.4 196.0 208.4 196.8 ;
      RECT  207.6 196.8 208.4 199.0 ;
      RECT  207.6 199.0 209.2 199.8 ;
      RECT  207.4 192.8 208.2 193.6 ;
      RECT  211.8 195.6 212.6 199.8 ;
      RECT  205.0 202.8 212.6 202.0 ;
      RECT  211.8 204.4 212.6 202.8 ;
      RECT  210.0 208.0 210.8 207.6 ;
      RECT  210.0 206.8 210.8 204.4 ;
      RECT  205.0 210.6 212.6 209.8 ;
      RECT  210.2 212.0 211.0 211.2 ;
      RECT  208.8 209.8 209.6 209.6 ;
      RECT  207.6 204.4 208.6 203.6 ;
      RECT  205.0 209.2 205.8 205.0 ;
      RECT  207.6 205.0 208.4 204.4 ;
      RECT  205.0 204.4 205.8 202.8 ;
      RECT  209.6 207.6 210.8 206.8 ;
      RECT  210.0 208.8 211.0 208.0 ;
      RECT  209.8 204.4 210.8 203.6 ;
      RECT  207.4 208.8 208.4 208.0 ;
      RECT  207.6 208.0 208.4 205.8 ;
      RECT  207.6 205.8 209.2 205.0 ;
      RECT  207.4 212.0 208.2 211.2 ;
      RECT  211.8 209.2 212.6 205.0 ;
      RECT  205.0 222.8 212.6 223.6 ;
      RECT  211.8 221.2 212.6 222.8 ;
      RECT  210.0 217.6 210.8 218.0 ;
      RECT  210.0 218.8 210.8 221.2 ;
      RECT  205.0 215.0 212.6 215.8 ;
      RECT  210.2 213.6 211.0 214.4 ;
      RECT  208.8 215.8 209.6 216.0 ;
      RECT  207.6 221.2 208.6 222.0 ;
      RECT  205.0 216.4 205.8 220.6 ;
      RECT  207.6 220.6 208.4 221.2 ;
      RECT  205.0 221.2 205.8 222.8 ;
      RECT  209.6 218.0 210.8 218.8 ;
      RECT  210.0 216.8 211.0 217.6 ;
      RECT  209.8 221.2 210.8 222.0 ;
      RECT  207.4 216.8 208.4 217.6 ;
      RECT  207.6 217.6 208.4 219.8 ;
      RECT  207.6 219.8 209.2 220.6 ;
      RECT  207.4 213.6 208.2 214.4 ;
      RECT  211.8 216.4 212.6 220.6 ;
      RECT  205.0 223.6 212.6 222.8 ;
      RECT  211.8 225.2 212.6 223.6 ;
      RECT  210.0 228.8 210.8 228.4 ;
      RECT  210.0 227.6 210.8 225.2 ;
      RECT  205.0 231.4 212.6 230.6 ;
      RECT  210.2 232.8 211.0 232.0 ;
      RECT  208.8 230.6 209.6 230.4 ;
      RECT  207.6 225.2 208.6 224.4 ;
      RECT  205.0 230.0 205.8 225.8 ;
      RECT  207.6 225.8 208.4 225.2 ;
      RECT  205.0 225.2 205.8 223.6 ;
      RECT  209.6 228.4 210.8 227.6 ;
      RECT  210.0 229.6 211.0 228.8 ;
      RECT  209.8 225.2 210.8 224.4 ;
      RECT  207.4 229.6 208.4 228.8 ;
      RECT  207.6 228.8 208.4 226.6 ;
      RECT  207.6 226.6 209.2 225.8 ;
      RECT  207.4 232.8 208.2 232.0 ;
      RECT  211.8 230.0 212.6 225.8 ;
      RECT  205.0 243.6 212.6 244.4 ;
      RECT  211.8 242.0 212.6 243.6 ;
      RECT  210.0 238.4 210.8 238.8 ;
      RECT  210.0 239.6 210.8 242.0 ;
      RECT  205.0 235.8 212.6 236.6 ;
      RECT  210.2 234.4 211.0 235.2 ;
      RECT  208.8 236.6 209.6 236.8 ;
      RECT  207.6 242.0 208.6 242.8 ;
      RECT  205.0 237.2 205.8 241.4 ;
      RECT  207.6 241.4 208.4 242.0 ;
      RECT  205.0 242.0 205.8 243.6 ;
      RECT  209.6 238.8 210.8 239.6 ;
      RECT  210.0 237.6 211.0 238.4 ;
      RECT  209.8 242.0 210.8 242.8 ;
      RECT  207.4 237.6 208.4 238.4 ;
      RECT  207.6 238.4 208.4 240.6 ;
      RECT  207.6 240.6 209.2 241.4 ;
      RECT  207.4 234.4 208.2 235.2 ;
      RECT  211.8 237.2 212.6 241.4 ;
      RECT  205.0 244.4 212.6 243.6 ;
      RECT  211.8 246.0 212.6 244.4 ;
      RECT  210.0 249.6 210.8 249.2 ;
      RECT  210.0 248.4 210.8 246.0 ;
      RECT  205.0 252.2 212.6 251.4 ;
      RECT  210.2 253.6 211.0 252.8 ;
      RECT  208.8 251.4 209.6 251.2 ;
      RECT  207.6 246.0 208.6 245.2 ;
      RECT  205.0 250.8 205.8 246.6 ;
      RECT  207.6 246.6 208.4 246.0 ;
      RECT  205.0 246.0 205.8 244.4 ;
      RECT  209.6 249.2 210.8 248.4 ;
      RECT  210.0 250.4 211.0 249.6 ;
      RECT  209.8 246.0 210.8 245.2 ;
      RECT  207.4 250.4 208.4 249.6 ;
      RECT  207.6 249.6 208.4 247.4 ;
      RECT  207.6 247.4 209.2 246.6 ;
      RECT  207.4 253.6 208.2 252.8 ;
      RECT  211.8 250.8 212.6 246.6 ;
      RECT  205.0 264.4 212.6 265.2 ;
      RECT  211.8 262.8 212.6 264.4 ;
      RECT  210.0 259.2 210.8 259.6 ;
      RECT  210.0 260.4 210.8 262.8 ;
      RECT  205.0 256.6 212.6 257.4 ;
      RECT  210.2 255.2 211.0 256.0 ;
      RECT  208.8 257.4 209.6 257.6 ;
      RECT  207.6 262.8 208.6 263.6 ;
      RECT  205.0 258.0 205.8 262.2 ;
      RECT  207.6 262.2 208.4 262.8 ;
      RECT  205.0 262.8 205.8 264.4 ;
      RECT  209.6 259.6 210.8 260.4 ;
      RECT  210.0 258.4 211.0 259.2 ;
      RECT  209.8 262.8 210.8 263.6 ;
      RECT  207.4 258.4 208.4 259.2 ;
      RECT  207.6 259.2 208.4 261.4 ;
      RECT  207.6 261.4 209.2 262.2 ;
      RECT  207.4 255.2 208.2 256.0 ;
      RECT  211.8 258.0 212.6 262.2 ;
      RECT  205.0 265.2 212.6 264.4 ;
      RECT  211.8 266.8 212.6 265.2 ;
      RECT  210.0 270.4 210.8 270.0 ;
      RECT  210.0 269.2 210.8 266.8 ;
      RECT  205.0 273.0 212.6 272.2 ;
      RECT  210.2 274.4 211.0 273.6 ;
      RECT  208.8 272.2 209.6 272.0 ;
      RECT  207.6 266.8 208.6 266.0 ;
      RECT  205.0 271.6 205.8 267.4 ;
      RECT  207.6 267.4 208.4 266.8 ;
      RECT  205.0 266.8 205.8 265.2 ;
      RECT  209.6 270.0 210.8 269.2 ;
      RECT  210.0 271.2 211.0 270.4 ;
      RECT  209.8 266.8 210.8 266.0 ;
      RECT  207.4 271.2 208.4 270.4 ;
      RECT  207.6 270.4 208.4 268.2 ;
      RECT  207.6 268.2 209.2 267.4 ;
      RECT  207.4 274.4 208.2 273.6 ;
      RECT  211.8 271.6 212.6 267.4 ;
      RECT  205.0 285.2 212.6 286.0 ;
      RECT  211.8 283.6 212.6 285.2 ;
      RECT  210.0 280.0 210.8 280.4 ;
      RECT  210.0 281.2 210.8 283.6 ;
      RECT  205.0 277.4 212.6 278.2 ;
      RECT  210.2 276.0 211.0 276.8 ;
      RECT  208.8 278.2 209.6 278.4 ;
      RECT  207.6 283.6 208.6 284.4 ;
      RECT  205.0 278.8 205.8 283.0 ;
      RECT  207.6 283.0 208.4 283.6 ;
      RECT  205.0 283.6 205.8 285.2 ;
      RECT  209.6 280.4 210.8 281.2 ;
      RECT  210.0 279.2 211.0 280.0 ;
      RECT  209.8 283.6 210.8 284.4 ;
      RECT  207.4 279.2 208.4 280.0 ;
      RECT  207.6 280.0 208.4 282.2 ;
      RECT  207.6 282.2 209.2 283.0 ;
      RECT  207.4 276.0 208.2 276.8 ;
      RECT  211.8 278.8 212.6 283.0 ;
      RECT  205.0 286.0 212.6 285.2 ;
      RECT  211.8 287.6 212.6 286.0 ;
      RECT  210.0 291.2 210.8 290.8 ;
      RECT  210.0 290.0 210.8 287.6 ;
      RECT  205.0 293.8 212.6 293.0 ;
      RECT  210.2 295.2 211.0 294.4 ;
      RECT  208.8 293.0 209.6 292.8 ;
      RECT  207.6 287.6 208.6 286.8 ;
      RECT  205.0 292.4 205.8 288.2 ;
      RECT  207.6 288.2 208.4 287.6 ;
      RECT  205.0 287.6 205.8 286.0 ;
      RECT  209.6 290.8 210.8 290.0 ;
      RECT  210.0 292.0 211.0 291.2 ;
      RECT  209.8 287.6 210.8 286.8 ;
      RECT  207.4 292.0 208.4 291.2 ;
      RECT  207.6 291.2 208.4 289.0 ;
      RECT  207.6 289.0 209.2 288.2 ;
      RECT  207.4 295.2 208.2 294.4 ;
      RECT  211.8 292.4 212.6 288.2 ;
      RECT  205.0 306.0 212.6 306.8 ;
      RECT  211.8 304.4 212.6 306.0 ;
      RECT  210.0 300.8 210.8 301.2 ;
      RECT  210.0 302.0 210.8 304.4 ;
      RECT  205.0 298.2 212.6 299.0 ;
      RECT  210.2 296.8 211.0 297.6 ;
      RECT  208.8 299.0 209.6 299.2 ;
      RECT  207.6 304.4 208.6 305.2 ;
      RECT  205.0 299.6 205.8 303.8 ;
      RECT  207.6 303.8 208.4 304.4 ;
      RECT  205.0 304.4 205.8 306.0 ;
      RECT  209.6 301.2 210.8 302.0 ;
      RECT  210.0 300.0 211.0 300.8 ;
      RECT  209.8 304.4 210.8 305.2 ;
      RECT  207.4 300.0 208.4 300.8 ;
      RECT  207.6 300.8 208.4 303.0 ;
      RECT  207.6 303.0 209.2 303.8 ;
      RECT  207.4 296.8 208.2 297.6 ;
      RECT  211.8 299.6 212.6 303.8 ;
      RECT  205.0 306.8 212.6 306.0 ;
      RECT  211.8 308.4 212.6 306.8 ;
      RECT  210.0 312.0 210.8 311.6 ;
      RECT  210.0 310.8 210.8 308.4 ;
      RECT  205.0 314.6 212.6 313.8 ;
      RECT  210.2 316.0 211.0 315.2 ;
      RECT  208.8 313.8 209.6 313.6 ;
      RECT  207.6 308.4 208.6 307.6 ;
      RECT  205.0 313.2 205.8 309.0 ;
      RECT  207.6 309.0 208.4 308.4 ;
      RECT  205.0 308.4 205.8 306.8 ;
      RECT  209.6 311.6 210.8 310.8 ;
      RECT  210.0 312.8 211.0 312.0 ;
      RECT  209.8 308.4 210.8 307.6 ;
      RECT  207.4 312.8 208.4 312.0 ;
      RECT  207.6 312.0 208.4 309.8 ;
      RECT  207.6 309.8 209.2 309.0 ;
      RECT  207.4 316.0 208.2 315.2 ;
      RECT  211.8 313.2 212.6 309.0 ;
      RECT  205.0 326.8 212.6 327.6 ;
      RECT  211.8 325.2 212.6 326.8 ;
      RECT  210.0 321.6 210.8 322.0 ;
      RECT  210.0 322.8 210.8 325.2 ;
      RECT  205.0 319.0 212.6 319.8 ;
      RECT  210.2 317.6 211.0 318.4 ;
      RECT  208.8 319.8 209.6 320.0 ;
      RECT  207.6 325.2 208.6 326.0 ;
      RECT  205.0 320.4 205.8 324.6 ;
      RECT  207.6 324.6 208.4 325.2 ;
      RECT  205.0 325.2 205.8 326.8 ;
      RECT  209.6 322.0 210.8 322.8 ;
      RECT  210.0 320.8 211.0 321.6 ;
      RECT  209.8 325.2 210.8 326.0 ;
      RECT  207.4 320.8 208.4 321.6 ;
      RECT  207.6 321.6 208.4 323.8 ;
      RECT  207.6 323.8 209.2 324.6 ;
      RECT  207.4 317.6 208.2 318.4 ;
      RECT  211.8 320.4 212.6 324.6 ;
      RECT  205.0 327.6 212.6 326.8 ;
      RECT  211.8 329.2 212.6 327.6 ;
      RECT  210.0 332.8 210.8 332.4 ;
      RECT  210.0 331.6 210.8 329.2 ;
      RECT  205.0 335.4 212.6 334.6 ;
      RECT  210.2 336.8 211.0 336.0 ;
      RECT  208.8 334.6 209.6 334.4 ;
      RECT  207.6 329.2 208.6 328.4 ;
      RECT  205.0 334.0 205.8 329.8 ;
      RECT  207.6 329.8 208.4 329.2 ;
      RECT  205.0 329.2 205.8 327.6 ;
      RECT  209.6 332.4 210.8 331.6 ;
      RECT  210.0 333.6 211.0 332.8 ;
      RECT  209.8 329.2 210.8 328.4 ;
      RECT  207.4 333.6 208.4 332.8 ;
      RECT  207.6 332.8 208.4 330.6 ;
      RECT  207.6 330.6 209.2 329.8 ;
      RECT  207.4 336.8 208.2 336.0 ;
      RECT  211.8 334.0 212.6 329.8 ;
      RECT  205.0 347.6 212.6 348.4 ;
      RECT  211.8 346.0 212.6 347.6 ;
      RECT  210.0 342.4 210.8 342.8 ;
      RECT  210.0 343.6 210.8 346.0 ;
      RECT  205.0 339.8 212.6 340.6 ;
      RECT  210.2 338.4 211.0 339.2 ;
      RECT  208.8 340.6 209.6 340.8 ;
      RECT  207.6 346.0 208.6 346.8 ;
      RECT  205.0 341.2 205.8 345.4 ;
      RECT  207.6 345.4 208.4 346.0 ;
      RECT  205.0 346.0 205.8 347.6 ;
      RECT  209.6 342.8 210.8 343.6 ;
      RECT  210.0 341.6 211.0 342.4 ;
      RECT  209.8 346.0 210.8 346.8 ;
      RECT  207.4 341.6 208.4 342.4 ;
      RECT  207.6 342.4 208.4 344.6 ;
      RECT  207.6 344.6 209.2 345.4 ;
      RECT  207.4 338.4 208.2 339.2 ;
      RECT  211.8 341.2 212.6 345.4 ;
      RECT  205.0 348.4 212.6 347.6 ;
      RECT  211.8 350.0 212.6 348.4 ;
      RECT  210.0 353.6 210.8 353.2 ;
      RECT  210.0 352.4 210.8 350.0 ;
      RECT  205.0 356.2 212.6 355.4 ;
      RECT  210.2 357.6 211.0 356.8 ;
      RECT  208.8 355.4 209.6 355.2 ;
      RECT  207.6 350.0 208.6 349.2 ;
      RECT  205.0 354.8 205.8 350.6 ;
      RECT  207.6 350.6 208.4 350.0 ;
      RECT  205.0 350.0 205.8 348.4 ;
      RECT  209.6 353.2 210.8 352.4 ;
      RECT  210.0 354.4 211.0 353.6 ;
      RECT  209.8 350.0 210.8 349.2 ;
      RECT  207.4 354.4 208.4 353.6 ;
      RECT  207.6 353.6 208.4 351.4 ;
      RECT  207.6 351.4 209.2 350.6 ;
      RECT  207.4 357.6 208.2 356.8 ;
      RECT  211.8 354.8 212.6 350.6 ;
      RECT  205.0 368.4 212.6 369.2 ;
      RECT  211.8 366.8 212.6 368.4 ;
      RECT  210.0 363.2 210.8 363.6 ;
      RECT  210.0 364.4 210.8 366.8 ;
      RECT  205.0 360.6 212.6 361.4 ;
      RECT  210.2 359.2 211.0 360.0 ;
      RECT  208.8 361.4 209.6 361.6 ;
      RECT  207.6 366.8 208.6 367.6 ;
      RECT  205.0 362.0 205.8 366.2 ;
      RECT  207.6 366.2 208.4 366.8 ;
      RECT  205.0 366.8 205.8 368.4 ;
      RECT  209.6 363.6 210.8 364.4 ;
      RECT  210.0 362.4 211.0 363.2 ;
      RECT  209.8 366.8 210.8 367.6 ;
      RECT  207.4 362.4 208.4 363.2 ;
      RECT  207.6 363.2 208.4 365.4 ;
      RECT  207.6 365.4 209.2 366.2 ;
      RECT  207.4 359.2 208.2 360.0 ;
      RECT  211.8 362.0 212.6 366.2 ;
      RECT  205.4 173.4 212.2 174.2 ;
      RECT  205.4 189.0 212.2 189.8 ;
      RECT  205.4 194.2 212.2 195.0 ;
      RECT  205.4 209.8 212.2 210.6 ;
      RECT  205.4 215.0 212.2 215.8 ;
      RECT  205.4 230.6 212.2 231.4 ;
      RECT  205.4 235.8 212.2 236.6 ;
      RECT  205.4 251.4 212.2 252.2 ;
      RECT  205.4 256.6 212.2 257.4 ;
      RECT  205.4 272.2 212.2 273.0 ;
      RECT  205.4 277.4 212.2 278.2 ;
      RECT  205.4 293.0 212.2 293.8 ;
      RECT  205.4 298.2 212.2 299.0 ;
      RECT  205.4 313.8 212.2 314.6 ;
      RECT  205.4 319.0 212.2 319.8 ;
      RECT  205.4 334.6 212.2 335.4 ;
      RECT  205.4 339.8 212.2 340.6 ;
      RECT  205.4 355.4 212.2 356.2 ;
      RECT  205.4 360.6 212.2 361.4 ;
      RECT  178.2 194.2 212.2 195.0 ;
      RECT  178.2 209.8 212.2 210.6 ;
      RECT  178.2 215.0 212.2 215.8 ;
      RECT  178.2 230.6 212.2 231.4 ;
      RECT  178.2 235.8 212.2 236.6 ;
      RECT  178.2 251.4 212.2 252.2 ;
      RECT  178.2 256.6 212.2 257.4 ;
      RECT  178.2 272.2 212.2 273.0 ;
      RECT  178.2 277.4 212.2 278.2 ;
      RECT  178.2 293.0 212.2 293.8 ;
      RECT  178.2 298.2 212.2 299.0 ;
      RECT  178.2 313.8 212.2 314.6 ;
      RECT  178.2 319.0 212.2 319.8 ;
      RECT  178.2 334.6 212.2 335.4 ;
      RECT  178.2 339.8 212.2 340.6 ;
      RECT  178.2 355.4 212.2 356.2 ;
      RECT  178.2 189.0 212.2 189.8 ;
      RECT  187.8 156.0 188.6 156.8 ;
      RECT  186.2 156.0 187.0 156.8 ;
      RECT  187.8 160.8 188.6 161.6 ;
      RECT  186.2 160.8 187.0 161.6 ;
      RECT  189.4 160.8 190.2 161.6 ;
      RECT  187.8 160.8 188.6 161.6 ;
      RECT  185.0 157.6 191.8 158.2 ;
      RECT  194.6 156.0 195.4 156.8 ;
      RECT  193.0 156.0 193.8 156.8 ;
      RECT  194.6 160.8 195.4 161.6 ;
      RECT  193.0 160.8 193.8 161.6 ;
      RECT  196.2 160.8 197.0 161.6 ;
      RECT  194.6 160.8 195.4 161.6 ;
      RECT  191.8 157.6 198.6 158.2 ;
      RECT  201.4 156.0 202.2 156.8 ;
      RECT  199.8 156.0 200.6 156.8 ;
      RECT  201.4 160.8 202.2 161.6 ;
      RECT  199.8 160.8 200.6 161.6 ;
      RECT  203.0 160.8 203.8 161.6 ;
      RECT  201.4 160.8 202.2 161.6 ;
      RECT  198.6 157.6 205.4 158.2 ;
      RECT  185.0 157.6 205.4 158.2 ;
      RECT  196.4 138.6 197.2 141.0 ;
      RECT  193.0 127.8 194.4 128.4 ;
      RECT  194.8 139.2 195.6 141.0 ;
      RECT  197.2 130.8 198.0 132.0 ;
      RECT  193.0 126.4 193.6 127.8 ;
      RECT  192.4 121.6 193.8 122.2 ;
      RECT  198.0 126.4 198.6 127.8 ;
      RECT  195.0 143.6 195.8 145.4 ;
      RECT  191.4 147.4 199.0 148.2 ;
      RECT  193.6 128.4 194.4 128.6 ;
      RECT  193.0 122.2 193.8 126.4 ;
      RECT  193.2 130.6 194.4 131.4 ;
      RECT  196.2 121.6 197.0 127.2 ;
      RECT  194.8 132.0 198.0 132.6 ;
      RECT  194.4 126.4 195.2 127.2 ;
      RECT  196.4 137.8 197.8 138.6 ;
      RECT  198.2 145.0 199.0 145.8 ;
      RECT  196.6 144.2 199.0 145.0 ;
      RECT  195.0 141.0 195.6 143.6 ;
      RECT  194.6 121.6 195.4 126.4 ;
      RECT  197.8 121.6 198.6 126.4 ;
      RECT  196.4 133.2 197.2 137.8 ;
      RECT  197.6 127.8 198.6 128.6 ;
      RECT  192.4 119.8 193.2 121.6 ;
      RECT  196.6 145.0 197.4 145.4 ;
      RECT  193.2 131.4 194.0 141.0 ;
      RECT  194.8 132.6 195.4 133.2 ;
      RECT  196.6 143.6 197.4 144.2 ;
      RECT  194.8 133.2 195.6 136.8 ;
      RECT  203.2 138.6 204.0 141.0 ;
      RECT  199.8 127.8 201.2 128.4 ;
      RECT  201.6 139.2 202.4 141.0 ;
      RECT  204.0 130.8 204.8 132.0 ;
      RECT  199.8 126.4 200.4 127.8 ;
      RECT  199.2 121.6 200.6 122.2 ;
      RECT  204.8 126.4 205.4 127.8 ;
      RECT  201.8 143.6 202.6 145.4 ;
      RECT  198.2 147.4 205.8 148.2 ;
      RECT  200.4 128.4 201.2 128.6 ;
      RECT  199.8 122.2 200.6 126.4 ;
      RECT  200.0 130.6 201.2 131.4 ;
      RECT  203.0 121.6 203.8 127.2 ;
      RECT  201.6 132.0 204.8 132.6 ;
      RECT  201.2 126.4 202.0 127.2 ;
      RECT  203.2 137.8 204.6 138.6 ;
      RECT  205.0 145.0 205.8 145.8 ;
      RECT  203.4 144.2 205.8 145.0 ;
      RECT  201.8 141.0 202.4 143.6 ;
      RECT  201.4 121.6 202.2 126.4 ;
      RECT  204.6 121.6 205.4 126.4 ;
      RECT  203.2 133.2 204.0 137.8 ;
      RECT  204.4 127.8 205.4 128.6 ;
      RECT  199.2 119.8 200.0 121.6 ;
      RECT  203.4 145.0 204.2 145.4 ;
      RECT  200.0 131.4 200.8 141.0 ;
      RECT  201.6 132.6 202.2 133.2 ;
      RECT  203.4 143.6 204.2 144.2 ;
      RECT  201.6 133.2 202.4 136.8 ;
      RECT  191.8 147.4 205.4 148.0 ;
      RECT  195.6 84.2 196.4 86.4 ;
      RECT  194.2 96.4 195.8 97.2 ;
      RECT  196.0 92.0 197.2 92.8 ;
      RECT  192.8 89.2 193.6 93.0 ;
      RECT  194.2 97.2 195.0 99.2 ;
      RECT  196.0 89.2 197.8 90.6 ;
      RECT  196.4 87.8 198.0 88.6 ;
      RECT  192.8 93.0 196.8 93.6 ;
      RECT  196.0 92.8 196.8 93.0 ;
      RECT  194.0 84.2 194.8 85.6 ;
      RECT  192.6 108.4 193.4 110.8 ;
      RECT  192.8 93.6 193.6 95.6 ;
      RECT  196.0 93.6 196.8 95.6 ;
      RECT  194.0 80.4 194.8 82.4 ;
      RECT  194.4 89.2 195.2 90.6 ;
      RECT  192.4 83.0 193.2 85.6 ;
      RECT  195.8 101.2 196.6 102.4 ;
      RECT  192.4 87.0 193.2 87.8 ;
      RECT  192.4 79.0 196.4 79.8 ;
      RECT  194.8 74.0 195.6 75.6 ;
      RECT  195.8 97.8 196.6 100.4 ;
      RECT  195.8 108.4 196.6 111.6 ;
      RECT  192.4 79.8 193.2 81.8 ;
      RECT  195.6 79.8 196.4 81.8 ;
      RECT  195.8 100.4 198.4 101.2 ;
      RECT  197.4 109.2 198.4 110.0 ;
      RECT  192.6 97.8 193.4 106.4 ;
      RECT  192.4 82.4 194.8 83.0 ;
      RECT  194.2 101.6 195.0 110.8 ;
      RECT  196.8 90.6 197.8 90.8 ;
      RECT  192.4 77.6 198.0 78.4 ;
      RECT  197.8 101.2 198.4 109.2 ;
      RECT  194.4 94.2 195.2 96.4 ;
      RECT  197.2 80.4 198.0 87.8 ;
      RECT  192.8 110.8 193.4 111.4 ;
      RECT  192.6 85.6 193.2 87.0 ;
      RECT  192.8 111.4 194.6 112.2 ;
      RECT  202.4 84.2 203.2 86.4 ;
      RECT  201.0 96.4 202.6 97.2 ;
      RECT  202.8 92.0 204.0 92.8 ;
      RECT  199.6 89.2 200.4 93.0 ;
      RECT  201.0 97.2 201.8 99.2 ;
      RECT  202.8 89.2 204.6 90.6 ;
      RECT  203.2 87.8 204.8 88.6 ;
      RECT  199.6 93.0 203.6 93.6 ;
      RECT  202.8 92.8 203.6 93.0 ;
      RECT  200.8 84.2 201.6 85.6 ;
      RECT  199.4 108.4 200.2 110.8 ;
      RECT  199.6 93.6 200.4 95.6 ;
      RECT  202.8 93.6 203.6 95.6 ;
      RECT  200.8 80.4 201.6 82.4 ;
      RECT  201.2 89.2 202.0 90.6 ;
      RECT  199.2 83.0 200.0 85.6 ;
      RECT  202.6 101.2 203.4 102.4 ;
      RECT  199.2 87.0 200.0 87.8 ;
      RECT  199.2 79.0 203.2 79.8 ;
      RECT  201.6 74.0 202.4 75.6 ;
      RECT  202.6 97.8 203.4 100.4 ;
      RECT  202.6 108.4 203.4 111.6 ;
      RECT  199.2 79.8 200.0 81.8 ;
      RECT  202.4 79.8 203.2 81.8 ;
      RECT  202.6 100.4 205.2 101.2 ;
      RECT  204.2 109.2 205.2 110.0 ;
      RECT  199.4 97.8 200.2 106.4 ;
      RECT  199.2 82.4 201.6 83.0 ;
      RECT  201.0 101.6 201.8 110.8 ;
      RECT  203.6 90.6 204.6 90.8 ;
      RECT  199.2 77.6 204.8 78.4 ;
      RECT  204.6 101.2 205.2 109.2 ;
      RECT  201.2 94.2 202.0 96.4 ;
      RECT  204.0 80.4 204.8 87.8 ;
      RECT  199.6 110.8 200.2 111.4 ;
      RECT  199.4 85.6 200.0 87.0 ;
      RECT  199.6 111.4 201.4 112.2 ;
      RECT  191.8 77.6 205.4 78.2 ;
      RECT  191.8 148.0 205.4 147.4 ;
      RECT  185.0 158.2 205.4 157.6 ;
      RECT  191.8 78.2 205.4 77.6 ;
      RECT  99.9 200.6 100.7 201.4 ;
      RECT  98.3 200.6 99.1 201.4 ;
      RECT  99.9 193.4 100.7 194.2 ;
      RECT  98.3 193.4 99.1 194.2 ;
      RECT  98.5 197.0 99.3 197.8 ;
      RECT  100.3 197.1 100.9 197.7 ;
      RECT  97.1 202.5 103.5 203.1 ;
      RECT  97.1 192.1 103.5 192.7 ;
      RECT  99.9 205.0 100.7 204.2 ;
      RECT  98.3 205.0 99.1 204.2 ;
      RECT  99.9 212.2 100.7 211.4 ;
      RECT  98.3 212.2 99.1 211.4 ;
      RECT  98.5 208.6 99.3 207.8 ;
      RECT  100.3 208.5 100.9 207.9 ;
      RECT  97.1 203.1 103.5 202.5 ;
      RECT  97.1 213.5 103.5 212.9 ;
      RECT  122.5 200.6 123.3 201.4 ;
      RECT  120.9 200.6 121.7 201.4 ;
      RECT  122.5 193.4 123.3 194.2 ;
      RECT  120.9 193.4 121.7 194.2 ;
      RECT  121.1 197.0 121.9 197.8 ;
      RECT  122.9 197.1 123.5 197.7 ;
      RECT  119.7 202.5 126.1 203.1 ;
      RECT  119.7 192.1 126.1 192.7 ;
      RECT  122.5 205.0 123.3 204.2 ;
      RECT  120.9 205.0 121.7 204.2 ;
      RECT  122.5 212.2 123.3 211.4 ;
      RECT  120.9 212.2 121.7 211.4 ;
      RECT  121.1 208.6 121.9 207.8 ;
      RECT  122.9 208.5 123.5 207.9 ;
      RECT  119.7 203.1 126.1 202.5 ;
      RECT  119.7 213.5 126.1 212.9 ;
      RECT  122.5 221.4 123.3 222.2 ;
      RECT  120.9 221.4 121.7 222.2 ;
      RECT  122.5 214.2 123.3 215.0 ;
      RECT  120.9 214.2 121.7 215.0 ;
      RECT  121.1 217.8 121.9 218.6 ;
      RECT  122.9 217.9 123.5 218.5 ;
      RECT  119.7 223.3 126.1 223.9 ;
      RECT  119.7 212.9 126.1 213.5 ;
      RECT  122.5 225.8 123.3 225.0 ;
      RECT  120.9 225.8 121.7 225.0 ;
      RECT  122.5 233.0 123.3 232.2 ;
      RECT  120.9 233.0 121.7 232.2 ;
      RECT  121.1 229.4 121.9 228.6 ;
      RECT  122.9 229.3 123.5 228.7 ;
      RECT  119.7 223.9 126.1 223.3 ;
      RECT  119.7 234.3 126.1 233.7 ;
      RECT  114.7 200.6 115.5 201.4 ;
      RECT  113.1 200.6 113.9 201.4 ;
      RECT  116.3 200.6 117.1 201.4 ;
      RECT  114.7 200.6 115.5 201.4 ;
      RECT  114.7 193.8 115.5 194.6 ;
      RECT  113.1 193.8 113.9 194.6 ;
      RECT  116.3 193.8 117.1 194.6 ;
      RECT  114.7 193.8 115.5 194.6 ;
      RECT  113.5 196.9 114.3 197.7 ;
      RECT  115.5 195.5 116.3 196.3 ;
      RECT  117.7 196.9 118.5 197.7 ;
      RECT  111.9 202.5 119.7 203.1 ;
      RECT  111.9 192.1 119.7 192.7 ;
      RECT  114.7 205.0 115.5 204.2 ;
      RECT  113.1 205.0 113.9 204.2 ;
      RECT  116.3 205.0 117.1 204.2 ;
      RECT  114.7 205.0 115.5 204.2 ;
      RECT  114.7 211.8 115.5 211.0 ;
      RECT  113.1 211.8 113.9 211.0 ;
      RECT  116.3 211.8 117.1 211.0 ;
      RECT  114.7 211.8 115.5 211.0 ;
      RECT  113.5 208.7 114.3 207.9 ;
      RECT  115.5 210.1 116.3 209.3 ;
      RECT  117.7 208.7 118.5 207.9 ;
      RECT  111.9 203.1 119.7 202.5 ;
      RECT  111.9 213.5 119.7 212.9 ;
      RECT  114.7 221.4 115.5 222.2 ;
      RECT  113.1 221.4 113.9 222.2 ;
      RECT  116.3 221.4 117.1 222.2 ;
      RECT  114.7 221.4 115.5 222.2 ;
      RECT  114.7 214.6 115.5 215.4 ;
      RECT  113.1 214.6 113.9 215.4 ;
      RECT  116.3 214.6 117.1 215.4 ;
      RECT  114.7 214.6 115.5 215.4 ;
      RECT  113.5 217.7 114.3 218.5 ;
      RECT  115.5 216.3 116.3 217.1 ;
      RECT  117.7 217.7 118.5 218.5 ;
      RECT  111.9 223.3 119.7 223.9 ;
      RECT  111.9 212.9 119.7 213.5 ;
      RECT  114.7 225.8 115.5 225.0 ;
      RECT  113.1 225.8 113.9 225.0 ;
      RECT  116.3 225.8 117.1 225.0 ;
      RECT  114.7 225.8 115.5 225.0 ;
      RECT  114.7 232.6 115.5 231.8 ;
      RECT  113.1 232.6 113.9 231.8 ;
      RECT  116.3 232.6 117.1 231.8 ;
      RECT  114.7 232.6 115.5 231.8 ;
      RECT  113.5 229.5 114.3 228.7 ;
      RECT  115.5 230.9 116.3 230.1 ;
      RECT  117.7 229.5 118.5 228.7 ;
      RECT  111.9 223.9 119.7 223.3 ;
      RECT  111.9 234.3 119.7 233.7 ;
      RECT  122.9 197.1 123.5 197.7 ;
      RECT  122.9 207.9 123.5 208.5 ;
      RECT  122.9 217.9 123.5 218.5 ;
      RECT  122.9 228.7 123.5 229.3 ;
      RECT  99.9 242.2 100.7 243.0 ;
      RECT  98.3 242.2 99.1 243.0 ;
      RECT  99.9 235.0 100.7 235.8 ;
      RECT  98.3 235.0 99.1 235.8 ;
      RECT  98.5 238.6 99.3 239.4 ;
      RECT  100.3 238.7 100.9 239.3 ;
      RECT  97.1 244.1 103.5 244.7 ;
      RECT  97.1 233.7 103.5 234.3 ;
      RECT  99.9 246.6 100.7 245.8 ;
      RECT  98.3 246.6 99.1 245.8 ;
      RECT  99.9 253.8 100.7 253.0 ;
      RECT  98.3 253.8 99.1 253.0 ;
      RECT  98.5 250.2 99.3 249.4 ;
      RECT  100.3 250.1 100.9 249.5 ;
      RECT  97.1 244.7 103.5 244.1 ;
      RECT  97.1 255.1 103.5 254.5 ;
      RECT  122.5 242.2 123.3 243.0 ;
      RECT  120.9 242.2 121.7 243.0 ;
      RECT  122.5 235.0 123.3 235.8 ;
      RECT  120.9 235.0 121.7 235.8 ;
      RECT  121.1 238.6 121.9 239.4 ;
      RECT  122.9 238.7 123.5 239.3 ;
      RECT  119.7 244.1 126.1 244.7 ;
      RECT  119.7 233.7 126.1 234.3 ;
      RECT  122.5 246.6 123.3 245.8 ;
      RECT  120.9 246.6 121.7 245.8 ;
      RECT  122.5 253.8 123.3 253.0 ;
      RECT  120.9 253.8 121.7 253.0 ;
      RECT  121.1 250.2 121.9 249.4 ;
      RECT  122.9 250.1 123.5 249.5 ;
      RECT  119.7 244.7 126.1 244.1 ;
      RECT  119.7 255.1 126.1 254.5 ;
      RECT  122.5 263.0 123.3 263.8 ;
      RECT  120.9 263.0 121.7 263.8 ;
      RECT  122.5 255.8 123.3 256.6 ;
      RECT  120.9 255.8 121.7 256.6 ;
      RECT  121.1 259.4 121.9 260.2 ;
      RECT  122.9 259.5 123.5 260.1 ;
      RECT  119.7 264.9 126.1 265.5 ;
      RECT  119.7 254.5 126.1 255.1 ;
      RECT  122.5 267.4 123.3 266.6 ;
      RECT  120.9 267.4 121.7 266.6 ;
      RECT  122.5 274.6 123.3 273.8 ;
      RECT  120.9 274.6 121.7 273.8 ;
      RECT  121.1 271.0 121.9 270.2 ;
      RECT  122.9 270.9 123.5 270.3 ;
      RECT  119.7 265.5 126.1 264.9 ;
      RECT  119.7 275.9 126.1 275.3 ;
      RECT  114.7 242.2 115.5 243.0 ;
      RECT  113.1 242.2 113.9 243.0 ;
      RECT  116.3 242.2 117.1 243.0 ;
      RECT  114.7 242.2 115.5 243.0 ;
      RECT  114.7 235.4 115.5 236.2 ;
      RECT  113.1 235.4 113.9 236.2 ;
      RECT  116.3 235.4 117.1 236.2 ;
      RECT  114.7 235.4 115.5 236.2 ;
      RECT  113.5 238.5 114.3 239.3 ;
      RECT  115.5 237.1 116.3 237.9 ;
      RECT  117.7 238.5 118.5 239.3 ;
      RECT  111.9 244.1 119.7 244.7 ;
      RECT  111.9 233.7 119.7 234.3 ;
      RECT  114.7 246.6 115.5 245.8 ;
      RECT  113.1 246.6 113.9 245.8 ;
      RECT  116.3 246.6 117.1 245.8 ;
      RECT  114.7 246.6 115.5 245.8 ;
      RECT  114.7 253.4 115.5 252.6 ;
      RECT  113.1 253.4 113.9 252.6 ;
      RECT  116.3 253.4 117.1 252.6 ;
      RECT  114.7 253.4 115.5 252.6 ;
      RECT  113.5 250.3 114.3 249.5 ;
      RECT  115.5 251.7 116.3 250.9 ;
      RECT  117.7 250.3 118.5 249.5 ;
      RECT  111.9 244.7 119.7 244.1 ;
      RECT  111.9 255.1 119.7 254.5 ;
      RECT  114.7 263.0 115.5 263.8 ;
      RECT  113.1 263.0 113.9 263.8 ;
      RECT  116.3 263.0 117.1 263.8 ;
      RECT  114.7 263.0 115.5 263.8 ;
      RECT  114.7 256.2 115.5 257.0 ;
      RECT  113.1 256.2 113.9 257.0 ;
      RECT  116.3 256.2 117.1 257.0 ;
      RECT  114.7 256.2 115.5 257.0 ;
      RECT  113.5 259.3 114.3 260.1 ;
      RECT  115.5 257.9 116.3 258.7 ;
      RECT  117.7 259.3 118.5 260.1 ;
      RECT  111.9 264.9 119.7 265.5 ;
      RECT  111.9 254.5 119.7 255.1 ;
      RECT  114.7 267.4 115.5 266.6 ;
      RECT  113.1 267.4 113.9 266.6 ;
      RECT  116.3 267.4 117.1 266.6 ;
      RECT  114.7 267.4 115.5 266.6 ;
      RECT  114.7 274.2 115.5 273.4 ;
      RECT  113.1 274.2 113.9 273.4 ;
      RECT  116.3 274.2 117.1 273.4 ;
      RECT  114.7 274.2 115.5 273.4 ;
      RECT  113.5 271.1 114.3 270.3 ;
      RECT  115.5 272.5 116.3 271.7 ;
      RECT  117.7 271.1 118.5 270.3 ;
      RECT  111.9 265.5 119.7 264.9 ;
      RECT  111.9 275.9 119.7 275.3 ;
      RECT  122.9 238.7 123.5 239.3 ;
      RECT  122.9 249.5 123.5 250.1 ;
      RECT  122.9 259.5 123.5 260.1 ;
      RECT  122.9 270.3 123.5 270.9 ;
      RECT  140.1 200.6 140.9 201.4 ;
      RECT  138.5 200.6 139.3 201.4 ;
      RECT  141.7 200.6 142.5 201.4 ;
      RECT  140.1 200.6 140.9 201.4 ;
      RECT  140.1 193.8 140.9 194.6 ;
      RECT  138.5 193.8 139.3 194.6 ;
      RECT  141.7 193.8 142.5 194.6 ;
      RECT  140.1 193.8 140.9 194.6 ;
      RECT  138.9 196.9 139.7 197.7 ;
      RECT  140.9 195.5 141.7 196.3 ;
      RECT  143.1 196.9 143.9 197.7 ;
      RECT  137.3 202.5 145.1 203.1 ;
      RECT  137.3 192.1 145.1 192.7 ;
      RECT  140.1 205.0 140.9 204.2 ;
      RECT  138.5 205.0 139.3 204.2 ;
      RECT  141.7 205.0 142.5 204.2 ;
      RECT  140.1 205.0 140.9 204.2 ;
      RECT  140.1 211.8 140.9 211.0 ;
      RECT  138.5 211.8 139.3 211.0 ;
      RECT  141.7 211.8 142.5 211.0 ;
      RECT  140.1 211.8 140.9 211.0 ;
      RECT  138.9 208.7 139.7 207.9 ;
      RECT  140.9 210.1 141.7 209.3 ;
      RECT  143.1 208.7 143.9 207.9 ;
      RECT  137.3 203.1 145.1 202.5 ;
      RECT  137.3 213.5 145.1 212.9 ;
      RECT  140.1 221.4 140.9 222.2 ;
      RECT  138.5 221.4 139.3 222.2 ;
      RECT  141.7 221.4 142.5 222.2 ;
      RECT  140.1 221.4 140.9 222.2 ;
      RECT  140.1 214.6 140.9 215.4 ;
      RECT  138.5 214.6 139.3 215.4 ;
      RECT  141.7 214.6 142.5 215.4 ;
      RECT  140.1 214.6 140.9 215.4 ;
      RECT  138.9 217.7 139.7 218.5 ;
      RECT  140.9 216.3 141.7 217.1 ;
      RECT  143.1 217.7 143.9 218.5 ;
      RECT  137.3 223.3 145.1 223.9 ;
      RECT  137.3 212.9 145.1 213.5 ;
      RECT  140.1 225.8 140.9 225.0 ;
      RECT  138.5 225.8 139.3 225.0 ;
      RECT  141.7 225.8 142.5 225.0 ;
      RECT  140.1 225.8 140.9 225.0 ;
      RECT  140.1 232.6 140.9 231.8 ;
      RECT  138.5 232.6 139.3 231.8 ;
      RECT  141.7 232.6 142.5 231.8 ;
      RECT  140.1 232.6 140.9 231.8 ;
      RECT  138.9 229.5 139.7 228.7 ;
      RECT  140.9 230.9 141.7 230.1 ;
      RECT  143.1 229.5 143.9 228.7 ;
      RECT  137.3 223.9 145.1 223.3 ;
      RECT  137.3 234.3 145.1 233.7 ;
      RECT  140.1 242.2 140.9 243.0 ;
      RECT  138.5 242.2 139.3 243.0 ;
      RECT  141.7 242.2 142.5 243.0 ;
      RECT  140.1 242.2 140.9 243.0 ;
      RECT  140.1 235.4 140.9 236.2 ;
      RECT  138.5 235.4 139.3 236.2 ;
      RECT  141.7 235.4 142.5 236.2 ;
      RECT  140.1 235.4 140.9 236.2 ;
      RECT  138.9 238.5 139.7 239.3 ;
      RECT  140.9 237.1 141.7 237.9 ;
      RECT  143.1 238.5 143.9 239.3 ;
      RECT  137.3 244.1 145.1 244.7 ;
      RECT  137.3 233.7 145.1 234.3 ;
      RECT  140.1 246.6 140.9 245.8 ;
      RECT  138.5 246.6 139.3 245.8 ;
      RECT  141.7 246.6 142.5 245.8 ;
      RECT  140.1 246.6 140.9 245.8 ;
      RECT  140.1 253.4 140.9 252.6 ;
      RECT  138.5 253.4 139.3 252.6 ;
      RECT  141.7 253.4 142.5 252.6 ;
      RECT  140.1 253.4 140.9 252.6 ;
      RECT  138.9 250.3 139.7 249.5 ;
      RECT  140.9 251.7 141.7 250.9 ;
      RECT  143.1 250.3 143.9 249.5 ;
      RECT  137.3 244.7 145.1 244.1 ;
      RECT  137.3 255.1 145.1 254.5 ;
      RECT  140.1 263.0 140.9 263.8 ;
      RECT  138.5 263.0 139.3 263.8 ;
      RECT  141.7 263.0 142.5 263.8 ;
      RECT  140.1 263.0 140.9 263.8 ;
      RECT  140.1 256.2 140.9 257.0 ;
      RECT  138.5 256.2 139.3 257.0 ;
      RECT  141.7 256.2 142.5 257.0 ;
      RECT  140.1 256.2 140.9 257.0 ;
      RECT  138.9 259.3 139.7 260.1 ;
      RECT  140.9 257.9 141.7 258.7 ;
      RECT  143.1 259.3 143.9 260.1 ;
      RECT  137.3 264.9 145.1 265.5 ;
      RECT  137.3 254.5 145.1 255.1 ;
      RECT  140.1 267.4 140.9 266.6 ;
      RECT  138.5 267.4 139.3 266.6 ;
      RECT  141.7 267.4 142.5 266.6 ;
      RECT  140.1 267.4 140.9 266.6 ;
      RECT  140.1 274.2 140.9 273.4 ;
      RECT  138.5 274.2 139.3 273.4 ;
      RECT  141.7 274.2 142.5 273.4 ;
      RECT  140.1 274.2 140.9 273.4 ;
      RECT  138.9 271.1 139.7 270.3 ;
      RECT  140.9 272.5 141.7 271.7 ;
      RECT  143.1 271.1 143.9 270.3 ;
      RECT  137.3 265.5 145.1 264.9 ;
      RECT  137.3 275.9 145.1 275.3 ;
      RECT  140.1 283.8 140.9 284.6 ;
      RECT  138.5 283.8 139.3 284.6 ;
      RECT  141.7 283.8 142.5 284.6 ;
      RECT  140.1 283.8 140.9 284.6 ;
      RECT  140.1 277.0 140.9 277.8 ;
      RECT  138.5 277.0 139.3 277.8 ;
      RECT  141.7 277.0 142.5 277.8 ;
      RECT  140.1 277.0 140.9 277.8 ;
      RECT  138.9 280.1 139.7 280.9 ;
      RECT  140.9 278.7 141.7 279.5 ;
      RECT  143.1 280.1 143.9 280.9 ;
      RECT  137.3 285.7 145.1 286.3 ;
      RECT  137.3 275.3 145.1 275.9 ;
      RECT  140.1 288.2 140.9 287.4 ;
      RECT  138.5 288.2 139.3 287.4 ;
      RECT  141.7 288.2 142.5 287.4 ;
      RECT  140.1 288.2 140.9 287.4 ;
      RECT  140.1 295.0 140.9 294.2 ;
      RECT  138.5 295.0 139.3 294.2 ;
      RECT  141.7 295.0 142.5 294.2 ;
      RECT  140.1 295.0 140.9 294.2 ;
      RECT  138.9 291.9 139.7 291.1 ;
      RECT  140.9 293.3 141.7 292.5 ;
      RECT  143.1 291.9 143.9 291.1 ;
      RECT  137.3 286.3 145.1 285.7 ;
      RECT  137.3 296.7 145.1 296.1 ;
      RECT  140.1 304.6 140.9 305.4 ;
      RECT  138.5 304.6 139.3 305.4 ;
      RECT  141.7 304.6 142.5 305.4 ;
      RECT  140.1 304.6 140.9 305.4 ;
      RECT  140.1 297.8 140.9 298.6 ;
      RECT  138.5 297.8 139.3 298.6 ;
      RECT  141.7 297.8 142.5 298.6 ;
      RECT  140.1 297.8 140.9 298.6 ;
      RECT  138.9 300.9 139.7 301.7 ;
      RECT  140.9 299.5 141.7 300.3 ;
      RECT  143.1 300.9 143.9 301.7 ;
      RECT  137.3 306.5 145.1 307.1 ;
      RECT  137.3 296.1 145.1 296.7 ;
      RECT  140.1 309.0 140.9 308.2 ;
      RECT  138.5 309.0 139.3 308.2 ;
      RECT  141.7 309.0 142.5 308.2 ;
      RECT  140.1 309.0 140.9 308.2 ;
      RECT  140.1 315.8 140.9 315.0 ;
      RECT  138.5 315.8 139.3 315.0 ;
      RECT  141.7 315.8 142.5 315.0 ;
      RECT  140.1 315.8 140.9 315.0 ;
      RECT  138.9 312.7 139.7 311.9 ;
      RECT  140.9 314.1 141.7 313.3 ;
      RECT  143.1 312.7 143.9 311.9 ;
      RECT  137.3 307.1 145.1 306.5 ;
      RECT  137.3 317.5 145.1 316.9 ;
      RECT  140.1 325.4 140.9 326.2 ;
      RECT  138.5 325.4 139.3 326.2 ;
      RECT  141.7 325.4 142.5 326.2 ;
      RECT  140.1 325.4 140.9 326.2 ;
      RECT  140.1 318.6 140.9 319.4 ;
      RECT  138.5 318.6 139.3 319.4 ;
      RECT  141.7 318.6 142.5 319.4 ;
      RECT  140.1 318.6 140.9 319.4 ;
      RECT  138.9 321.7 139.7 322.5 ;
      RECT  140.9 320.3 141.7 321.1 ;
      RECT  143.1 321.7 143.9 322.5 ;
      RECT  137.3 327.3 145.1 327.9 ;
      RECT  137.3 316.9 145.1 317.5 ;
      RECT  140.1 329.8 140.9 329.0 ;
      RECT  138.5 329.8 139.3 329.0 ;
      RECT  141.7 329.8 142.5 329.0 ;
      RECT  140.1 329.8 140.9 329.0 ;
      RECT  140.1 336.6 140.9 335.8 ;
      RECT  138.5 336.6 139.3 335.8 ;
      RECT  141.7 336.6 142.5 335.8 ;
      RECT  140.1 336.6 140.9 335.8 ;
      RECT  138.9 333.5 139.7 332.7 ;
      RECT  140.9 334.9 141.7 334.1 ;
      RECT  143.1 333.5 143.9 332.7 ;
      RECT  137.3 327.9 145.1 327.3 ;
      RECT  137.3 338.3 145.1 337.7 ;
      RECT  140.1 346.2 140.9 347.0 ;
      RECT  138.5 346.2 139.3 347.0 ;
      RECT  141.7 346.2 142.5 347.0 ;
      RECT  140.1 346.2 140.9 347.0 ;
      RECT  140.1 339.4 140.9 340.2 ;
      RECT  138.5 339.4 139.3 340.2 ;
      RECT  141.7 339.4 142.5 340.2 ;
      RECT  140.1 339.4 140.9 340.2 ;
      RECT  138.9 342.5 139.7 343.3 ;
      RECT  140.9 341.1 141.7 341.9 ;
      RECT  143.1 342.5 143.9 343.3 ;
      RECT  137.3 348.1 145.1 348.7 ;
      RECT  137.3 337.7 145.1 338.3 ;
      RECT  140.1 350.6 140.9 349.8 ;
      RECT  138.5 350.6 139.3 349.8 ;
      RECT  141.7 350.6 142.5 349.8 ;
      RECT  140.1 350.6 140.9 349.8 ;
      RECT  140.1 357.4 140.9 356.6 ;
      RECT  138.5 357.4 139.3 356.6 ;
      RECT  141.7 357.4 142.5 356.6 ;
      RECT  140.1 357.4 140.9 356.6 ;
      RECT  138.9 354.3 139.7 353.5 ;
      RECT  140.9 355.7 141.7 354.9 ;
      RECT  143.1 354.3 143.9 353.5 ;
      RECT  137.3 348.7 145.1 348.1 ;
      RECT  137.3 359.1 145.1 358.5 ;
      RECT  147.9 200.6 148.7 201.4 ;
      RECT  146.3 200.6 147.1 201.4 ;
      RECT  147.9 193.4 148.7 194.2 ;
      RECT  146.3 193.4 147.1 194.2 ;
      RECT  146.5 197.0 147.3 197.8 ;
      RECT  148.3 197.1 148.9 197.7 ;
      RECT  145.1 202.5 151.5 203.1 ;
      RECT  145.1 192.1 151.5 192.7 ;
      RECT  147.9 205.0 148.7 204.2 ;
      RECT  146.3 205.0 147.1 204.2 ;
      RECT  147.9 212.2 148.7 211.4 ;
      RECT  146.3 212.2 147.1 211.4 ;
      RECT  146.5 208.6 147.3 207.8 ;
      RECT  148.3 208.5 148.9 207.9 ;
      RECT  145.1 203.1 151.5 202.5 ;
      RECT  145.1 213.5 151.5 212.9 ;
      RECT  147.9 221.4 148.7 222.2 ;
      RECT  146.3 221.4 147.1 222.2 ;
      RECT  147.9 214.2 148.7 215.0 ;
      RECT  146.3 214.2 147.1 215.0 ;
      RECT  146.5 217.8 147.3 218.6 ;
      RECT  148.3 217.9 148.9 218.5 ;
      RECT  145.1 223.3 151.5 223.9 ;
      RECT  145.1 212.9 151.5 213.5 ;
      RECT  147.9 225.8 148.7 225.0 ;
      RECT  146.3 225.8 147.1 225.0 ;
      RECT  147.9 233.0 148.7 232.2 ;
      RECT  146.3 233.0 147.1 232.2 ;
      RECT  146.5 229.4 147.3 228.6 ;
      RECT  148.3 229.3 148.9 228.7 ;
      RECT  145.1 223.9 151.5 223.3 ;
      RECT  145.1 234.3 151.5 233.7 ;
      RECT  147.9 242.2 148.7 243.0 ;
      RECT  146.3 242.2 147.1 243.0 ;
      RECT  147.9 235.0 148.7 235.8 ;
      RECT  146.3 235.0 147.1 235.8 ;
      RECT  146.5 238.6 147.3 239.4 ;
      RECT  148.3 238.7 148.9 239.3 ;
      RECT  145.1 244.1 151.5 244.7 ;
      RECT  145.1 233.7 151.5 234.3 ;
      RECT  147.9 246.6 148.7 245.8 ;
      RECT  146.3 246.6 147.1 245.8 ;
      RECT  147.9 253.8 148.7 253.0 ;
      RECT  146.3 253.8 147.1 253.0 ;
      RECT  146.5 250.2 147.3 249.4 ;
      RECT  148.3 250.1 148.9 249.5 ;
      RECT  145.1 244.7 151.5 244.1 ;
      RECT  145.1 255.1 151.5 254.5 ;
      RECT  147.9 263.0 148.7 263.8 ;
      RECT  146.3 263.0 147.1 263.8 ;
      RECT  147.9 255.8 148.7 256.6 ;
      RECT  146.3 255.8 147.1 256.6 ;
      RECT  146.5 259.4 147.3 260.2 ;
      RECT  148.3 259.5 148.9 260.1 ;
      RECT  145.1 264.9 151.5 265.5 ;
      RECT  145.1 254.5 151.5 255.1 ;
      RECT  147.9 267.4 148.7 266.6 ;
      RECT  146.3 267.4 147.1 266.6 ;
      RECT  147.9 274.6 148.7 273.8 ;
      RECT  146.3 274.6 147.1 273.8 ;
      RECT  146.5 271.0 147.3 270.2 ;
      RECT  148.3 270.9 148.9 270.3 ;
      RECT  145.1 265.5 151.5 264.9 ;
      RECT  145.1 275.9 151.5 275.3 ;
      RECT  147.9 283.8 148.7 284.6 ;
      RECT  146.3 283.8 147.1 284.6 ;
      RECT  147.9 276.6 148.7 277.4 ;
      RECT  146.3 276.6 147.1 277.4 ;
      RECT  146.5 280.2 147.3 281.0 ;
      RECT  148.3 280.3 148.9 280.9 ;
      RECT  145.1 285.7 151.5 286.3 ;
      RECT  145.1 275.3 151.5 275.9 ;
      RECT  147.9 288.2 148.7 287.4 ;
      RECT  146.3 288.2 147.1 287.4 ;
      RECT  147.9 295.4 148.7 294.6 ;
      RECT  146.3 295.4 147.1 294.6 ;
      RECT  146.5 291.8 147.3 291.0 ;
      RECT  148.3 291.7 148.9 291.1 ;
      RECT  145.1 286.3 151.5 285.7 ;
      RECT  145.1 296.7 151.5 296.1 ;
      RECT  147.9 304.6 148.7 305.4 ;
      RECT  146.3 304.6 147.1 305.4 ;
      RECT  147.9 297.4 148.7 298.2 ;
      RECT  146.3 297.4 147.1 298.2 ;
      RECT  146.5 301.0 147.3 301.8 ;
      RECT  148.3 301.1 148.9 301.7 ;
      RECT  145.1 306.5 151.5 307.1 ;
      RECT  145.1 296.1 151.5 296.7 ;
      RECT  147.9 309.0 148.7 308.2 ;
      RECT  146.3 309.0 147.1 308.2 ;
      RECT  147.9 316.2 148.7 315.4 ;
      RECT  146.3 316.2 147.1 315.4 ;
      RECT  146.5 312.6 147.3 311.8 ;
      RECT  148.3 312.5 148.9 311.9 ;
      RECT  145.1 307.1 151.5 306.5 ;
      RECT  145.1 317.5 151.5 316.9 ;
      RECT  147.9 325.4 148.7 326.2 ;
      RECT  146.3 325.4 147.1 326.2 ;
      RECT  147.9 318.2 148.7 319.0 ;
      RECT  146.3 318.2 147.1 319.0 ;
      RECT  146.5 321.8 147.3 322.6 ;
      RECT  148.3 321.9 148.9 322.5 ;
      RECT  145.1 327.3 151.5 327.9 ;
      RECT  145.1 316.9 151.5 317.5 ;
      RECT  147.9 329.8 148.7 329.0 ;
      RECT  146.3 329.8 147.1 329.0 ;
      RECT  147.9 337.0 148.7 336.2 ;
      RECT  146.3 337.0 147.1 336.2 ;
      RECT  146.5 333.4 147.3 332.6 ;
      RECT  148.3 333.3 148.9 332.7 ;
      RECT  145.1 327.9 151.5 327.3 ;
      RECT  145.1 338.3 151.5 337.7 ;
      RECT  147.9 346.2 148.7 347.0 ;
      RECT  146.3 346.2 147.1 347.0 ;
      RECT  147.9 339.0 148.7 339.8 ;
      RECT  146.3 339.0 147.1 339.8 ;
      RECT  146.5 342.6 147.3 343.4 ;
      RECT  148.3 342.7 148.9 343.3 ;
      RECT  145.1 348.1 151.5 348.7 ;
      RECT  145.1 337.7 151.5 338.3 ;
      RECT  147.9 350.6 148.7 349.8 ;
      RECT  146.3 350.6 147.1 349.8 ;
      RECT  147.9 357.8 148.7 357.0 ;
      RECT  146.3 357.8 147.1 357.0 ;
      RECT  146.5 354.2 147.3 353.4 ;
      RECT  148.3 354.1 148.9 353.5 ;
      RECT  145.1 348.7 151.5 348.1 ;
      RECT  145.1 359.1 151.5 358.5 ;
      RECT  148.3 197.1 148.9 197.7 ;
      RECT  148.3 207.9 148.9 208.5 ;
      RECT  148.3 217.9 148.9 218.5 ;
      RECT  148.3 228.7 148.9 229.3 ;
      RECT  148.3 238.7 148.9 239.3 ;
      RECT  148.3 249.5 148.9 250.1 ;
      RECT  148.3 259.5 148.9 260.1 ;
      RECT  148.3 270.3 148.9 270.9 ;
      RECT  148.3 280.3 148.9 280.9 ;
      RECT  148.3 291.1 148.9 291.7 ;
      RECT  148.3 301.1 148.9 301.7 ;
      RECT  148.3 311.9 148.9 312.5 ;
      RECT  148.3 321.9 148.9 322.5 ;
      RECT  148.3 332.7 148.9 333.3 ;
      RECT  148.3 342.7 148.9 343.3 ;
      RECT  148.3 353.5 148.9 354.1 ;
      RECT  160.9 200.6 161.7 201.4 ;
      RECT  159.3 200.6 160.1 201.4 ;
      RECT  162.5 200.6 163.3 201.4 ;
      RECT  160.9 200.6 161.7 201.4 ;
      RECT  160.9 193.8 161.7 194.6 ;
      RECT  159.3 193.8 160.1 194.6 ;
      RECT  162.5 193.8 163.3 194.6 ;
      RECT  160.9 193.8 161.7 194.6 ;
      RECT  159.7 196.9 160.5 197.7 ;
      RECT  161.7 195.5 162.5 196.3 ;
      RECT  163.9 196.9 164.7 197.7 ;
      RECT  158.1 202.5 165.9 203.1 ;
      RECT  158.1 192.1 165.9 192.7 ;
      RECT  168.7 200.6 169.5 201.4 ;
      RECT  167.1 200.6 167.9 201.4 ;
      RECT  168.7 193.4 169.5 194.2 ;
      RECT  167.1 193.4 167.9 194.2 ;
      RECT  167.3 197.0 168.1 197.8 ;
      RECT  169.1 197.1 169.7 197.7 ;
      RECT  165.9 202.5 172.3 203.1 ;
      RECT  165.9 192.1 172.3 192.7 ;
      RECT  167.3 197.0 168.1 197.8 ;
      RECT  169.1 197.1 169.7 197.7 ;
      RECT  165.9 202.5 166.5 203.1 ;
      RECT  165.9 192.1 166.5 192.7 ;
      RECT  160.9 205.0 161.7 204.2 ;
      RECT  159.3 205.0 160.1 204.2 ;
      RECT  162.5 205.0 163.3 204.2 ;
      RECT  160.9 205.0 161.7 204.2 ;
      RECT  160.9 211.8 161.7 211.0 ;
      RECT  159.3 211.8 160.1 211.0 ;
      RECT  162.5 211.8 163.3 211.0 ;
      RECT  160.9 211.8 161.7 211.0 ;
      RECT  159.7 208.7 160.5 207.9 ;
      RECT  161.7 210.1 162.5 209.3 ;
      RECT  163.9 208.7 164.7 207.9 ;
      RECT  158.1 203.1 165.9 202.5 ;
      RECT  158.1 213.5 165.9 212.9 ;
      RECT  168.7 205.0 169.5 204.2 ;
      RECT  167.1 205.0 167.9 204.2 ;
      RECT  168.7 212.2 169.5 211.4 ;
      RECT  167.1 212.2 167.9 211.4 ;
      RECT  167.3 208.6 168.1 207.8 ;
      RECT  169.1 208.5 169.7 207.9 ;
      RECT  165.9 203.1 172.3 202.5 ;
      RECT  165.9 213.5 172.3 212.9 ;
      RECT  167.3 208.6 168.1 207.8 ;
      RECT  169.1 208.5 169.7 207.9 ;
      RECT  165.9 203.1 166.5 202.5 ;
      RECT  165.9 213.5 166.5 212.9 ;
      RECT  160.9 221.4 161.7 222.2 ;
      RECT  159.3 221.4 160.1 222.2 ;
      RECT  162.5 221.4 163.3 222.2 ;
      RECT  160.9 221.4 161.7 222.2 ;
      RECT  160.9 214.6 161.7 215.4 ;
      RECT  159.3 214.6 160.1 215.4 ;
      RECT  162.5 214.6 163.3 215.4 ;
      RECT  160.9 214.6 161.7 215.4 ;
      RECT  159.7 217.7 160.5 218.5 ;
      RECT  161.7 216.3 162.5 217.1 ;
      RECT  163.9 217.7 164.7 218.5 ;
      RECT  158.1 223.3 165.9 223.9 ;
      RECT  158.1 212.9 165.9 213.5 ;
      RECT  168.7 221.4 169.5 222.2 ;
      RECT  167.1 221.4 167.9 222.2 ;
      RECT  168.7 214.2 169.5 215.0 ;
      RECT  167.1 214.2 167.9 215.0 ;
      RECT  167.3 217.8 168.1 218.6 ;
      RECT  169.1 217.9 169.7 218.5 ;
      RECT  165.9 223.3 172.3 223.9 ;
      RECT  165.9 212.9 172.3 213.5 ;
      RECT  167.3 217.8 168.1 218.6 ;
      RECT  169.1 217.9 169.7 218.5 ;
      RECT  165.9 223.3 166.5 223.9 ;
      RECT  165.9 212.9 166.5 213.5 ;
      RECT  160.9 225.8 161.7 225.0 ;
      RECT  159.3 225.8 160.1 225.0 ;
      RECT  162.5 225.8 163.3 225.0 ;
      RECT  160.9 225.8 161.7 225.0 ;
      RECT  160.9 232.6 161.7 231.8 ;
      RECT  159.3 232.6 160.1 231.8 ;
      RECT  162.5 232.6 163.3 231.8 ;
      RECT  160.9 232.6 161.7 231.8 ;
      RECT  159.7 229.5 160.5 228.7 ;
      RECT  161.7 230.9 162.5 230.1 ;
      RECT  163.9 229.5 164.7 228.7 ;
      RECT  158.1 223.9 165.9 223.3 ;
      RECT  158.1 234.3 165.9 233.7 ;
      RECT  168.7 225.8 169.5 225.0 ;
      RECT  167.1 225.8 167.9 225.0 ;
      RECT  168.7 233.0 169.5 232.2 ;
      RECT  167.1 233.0 167.9 232.2 ;
      RECT  167.3 229.4 168.1 228.6 ;
      RECT  169.1 229.3 169.7 228.7 ;
      RECT  165.9 223.9 172.3 223.3 ;
      RECT  165.9 234.3 172.3 233.7 ;
      RECT  167.3 229.4 168.1 228.6 ;
      RECT  169.1 229.3 169.7 228.7 ;
      RECT  165.9 223.9 166.5 223.3 ;
      RECT  165.9 234.3 166.5 233.7 ;
      RECT  160.9 242.2 161.7 243.0 ;
      RECT  159.3 242.2 160.1 243.0 ;
      RECT  162.5 242.2 163.3 243.0 ;
      RECT  160.9 242.2 161.7 243.0 ;
      RECT  160.9 235.4 161.7 236.2 ;
      RECT  159.3 235.4 160.1 236.2 ;
      RECT  162.5 235.4 163.3 236.2 ;
      RECT  160.9 235.4 161.7 236.2 ;
      RECT  159.7 238.5 160.5 239.3 ;
      RECT  161.7 237.1 162.5 237.9 ;
      RECT  163.9 238.5 164.7 239.3 ;
      RECT  158.1 244.1 165.9 244.7 ;
      RECT  158.1 233.7 165.9 234.3 ;
      RECT  168.7 242.2 169.5 243.0 ;
      RECT  167.1 242.2 167.9 243.0 ;
      RECT  168.7 235.0 169.5 235.8 ;
      RECT  167.1 235.0 167.9 235.8 ;
      RECT  167.3 238.6 168.1 239.4 ;
      RECT  169.1 238.7 169.7 239.3 ;
      RECT  165.9 244.1 172.3 244.7 ;
      RECT  165.9 233.7 172.3 234.3 ;
      RECT  167.3 238.6 168.1 239.4 ;
      RECT  169.1 238.7 169.7 239.3 ;
      RECT  165.9 244.1 166.5 244.7 ;
      RECT  165.9 233.7 166.5 234.3 ;
      RECT  160.9 246.6 161.7 245.8 ;
      RECT  159.3 246.6 160.1 245.8 ;
      RECT  162.5 246.6 163.3 245.8 ;
      RECT  160.9 246.6 161.7 245.8 ;
      RECT  160.9 253.4 161.7 252.6 ;
      RECT  159.3 253.4 160.1 252.6 ;
      RECT  162.5 253.4 163.3 252.6 ;
      RECT  160.9 253.4 161.7 252.6 ;
      RECT  159.7 250.3 160.5 249.5 ;
      RECT  161.7 251.7 162.5 250.9 ;
      RECT  163.9 250.3 164.7 249.5 ;
      RECT  158.1 244.7 165.9 244.1 ;
      RECT  158.1 255.1 165.9 254.5 ;
      RECT  168.7 246.6 169.5 245.8 ;
      RECT  167.1 246.6 167.9 245.8 ;
      RECT  168.7 253.8 169.5 253.0 ;
      RECT  167.1 253.8 167.9 253.0 ;
      RECT  167.3 250.2 168.1 249.4 ;
      RECT  169.1 250.1 169.7 249.5 ;
      RECT  165.9 244.7 172.3 244.1 ;
      RECT  165.9 255.1 172.3 254.5 ;
      RECT  167.3 250.2 168.1 249.4 ;
      RECT  169.1 250.1 169.7 249.5 ;
      RECT  165.9 244.7 166.5 244.1 ;
      RECT  165.9 255.1 166.5 254.5 ;
      RECT  160.9 263.0 161.7 263.8 ;
      RECT  159.3 263.0 160.1 263.8 ;
      RECT  162.5 263.0 163.3 263.8 ;
      RECT  160.9 263.0 161.7 263.8 ;
      RECT  160.9 256.2 161.7 257.0 ;
      RECT  159.3 256.2 160.1 257.0 ;
      RECT  162.5 256.2 163.3 257.0 ;
      RECT  160.9 256.2 161.7 257.0 ;
      RECT  159.7 259.3 160.5 260.1 ;
      RECT  161.7 257.9 162.5 258.7 ;
      RECT  163.9 259.3 164.7 260.1 ;
      RECT  158.1 264.9 165.9 265.5 ;
      RECT  158.1 254.5 165.9 255.1 ;
      RECT  168.7 263.0 169.5 263.8 ;
      RECT  167.1 263.0 167.9 263.8 ;
      RECT  168.7 255.8 169.5 256.6 ;
      RECT  167.1 255.8 167.9 256.6 ;
      RECT  167.3 259.4 168.1 260.2 ;
      RECT  169.1 259.5 169.7 260.1 ;
      RECT  165.9 264.9 172.3 265.5 ;
      RECT  165.9 254.5 172.3 255.1 ;
      RECT  167.3 259.4 168.1 260.2 ;
      RECT  169.1 259.5 169.7 260.1 ;
      RECT  165.9 264.9 166.5 265.5 ;
      RECT  165.9 254.5 166.5 255.1 ;
      RECT  160.9 267.4 161.7 266.6 ;
      RECT  159.3 267.4 160.1 266.6 ;
      RECT  162.5 267.4 163.3 266.6 ;
      RECT  160.9 267.4 161.7 266.6 ;
      RECT  160.9 274.2 161.7 273.4 ;
      RECT  159.3 274.2 160.1 273.4 ;
      RECT  162.5 274.2 163.3 273.4 ;
      RECT  160.9 274.2 161.7 273.4 ;
      RECT  159.7 271.1 160.5 270.3 ;
      RECT  161.7 272.5 162.5 271.7 ;
      RECT  163.9 271.1 164.7 270.3 ;
      RECT  158.1 265.5 165.9 264.9 ;
      RECT  158.1 275.9 165.9 275.3 ;
      RECT  168.7 267.4 169.5 266.6 ;
      RECT  167.1 267.4 167.9 266.6 ;
      RECT  168.7 274.6 169.5 273.8 ;
      RECT  167.1 274.6 167.9 273.8 ;
      RECT  167.3 271.0 168.1 270.2 ;
      RECT  169.1 270.9 169.7 270.3 ;
      RECT  165.9 265.5 172.3 264.9 ;
      RECT  165.9 275.9 172.3 275.3 ;
      RECT  167.3 271.0 168.1 270.2 ;
      RECT  169.1 270.9 169.7 270.3 ;
      RECT  165.9 265.5 166.5 264.9 ;
      RECT  165.9 275.9 166.5 275.3 ;
      RECT  160.9 283.8 161.7 284.6 ;
      RECT  159.3 283.8 160.1 284.6 ;
      RECT  162.5 283.8 163.3 284.6 ;
      RECT  160.9 283.8 161.7 284.6 ;
      RECT  160.9 277.0 161.7 277.8 ;
      RECT  159.3 277.0 160.1 277.8 ;
      RECT  162.5 277.0 163.3 277.8 ;
      RECT  160.9 277.0 161.7 277.8 ;
      RECT  159.7 280.1 160.5 280.9 ;
      RECT  161.7 278.7 162.5 279.5 ;
      RECT  163.9 280.1 164.7 280.9 ;
      RECT  158.1 285.7 165.9 286.3 ;
      RECT  158.1 275.3 165.9 275.9 ;
      RECT  168.7 283.8 169.5 284.6 ;
      RECT  167.1 283.8 167.9 284.6 ;
      RECT  168.7 276.6 169.5 277.4 ;
      RECT  167.1 276.6 167.9 277.4 ;
      RECT  167.3 280.2 168.1 281.0 ;
      RECT  169.1 280.3 169.7 280.9 ;
      RECT  165.9 285.7 172.3 286.3 ;
      RECT  165.9 275.3 172.3 275.9 ;
      RECT  167.3 280.2 168.1 281.0 ;
      RECT  169.1 280.3 169.7 280.9 ;
      RECT  165.9 285.7 166.5 286.3 ;
      RECT  165.9 275.3 166.5 275.9 ;
      RECT  160.9 288.2 161.7 287.4 ;
      RECT  159.3 288.2 160.1 287.4 ;
      RECT  162.5 288.2 163.3 287.4 ;
      RECT  160.9 288.2 161.7 287.4 ;
      RECT  160.9 295.0 161.7 294.2 ;
      RECT  159.3 295.0 160.1 294.2 ;
      RECT  162.5 295.0 163.3 294.2 ;
      RECT  160.9 295.0 161.7 294.2 ;
      RECT  159.7 291.9 160.5 291.1 ;
      RECT  161.7 293.3 162.5 292.5 ;
      RECT  163.9 291.9 164.7 291.1 ;
      RECT  158.1 286.3 165.9 285.7 ;
      RECT  158.1 296.7 165.9 296.1 ;
      RECT  168.7 288.2 169.5 287.4 ;
      RECT  167.1 288.2 167.9 287.4 ;
      RECT  168.7 295.4 169.5 294.6 ;
      RECT  167.1 295.4 167.9 294.6 ;
      RECT  167.3 291.8 168.1 291.0 ;
      RECT  169.1 291.7 169.7 291.1 ;
      RECT  165.9 286.3 172.3 285.7 ;
      RECT  165.9 296.7 172.3 296.1 ;
      RECT  167.3 291.8 168.1 291.0 ;
      RECT  169.1 291.7 169.7 291.1 ;
      RECT  165.9 286.3 166.5 285.7 ;
      RECT  165.9 296.7 166.5 296.1 ;
      RECT  160.9 304.6 161.7 305.4 ;
      RECT  159.3 304.6 160.1 305.4 ;
      RECT  162.5 304.6 163.3 305.4 ;
      RECT  160.9 304.6 161.7 305.4 ;
      RECT  160.9 297.8 161.7 298.6 ;
      RECT  159.3 297.8 160.1 298.6 ;
      RECT  162.5 297.8 163.3 298.6 ;
      RECT  160.9 297.8 161.7 298.6 ;
      RECT  159.7 300.9 160.5 301.7 ;
      RECT  161.7 299.5 162.5 300.3 ;
      RECT  163.9 300.9 164.7 301.7 ;
      RECT  158.1 306.5 165.9 307.1 ;
      RECT  158.1 296.1 165.9 296.7 ;
      RECT  168.7 304.6 169.5 305.4 ;
      RECT  167.1 304.6 167.9 305.4 ;
      RECT  168.7 297.4 169.5 298.2 ;
      RECT  167.1 297.4 167.9 298.2 ;
      RECT  167.3 301.0 168.1 301.8 ;
      RECT  169.1 301.1 169.7 301.7 ;
      RECT  165.9 306.5 172.3 307.1 ;
      RECT  165.9 296.1 172.3 296.7 ;
      RECT  167.3 301.0 168.1 301.8 ;
      RECT  169.1 301.1 169.7 301.7 ;
      RECT  165.9 306.5 166.5 307.1 ;
      RECT  165.9 296.1 166.5 296.7 ;
      RECT  160.9 309.0 161.7 308.2 ;
      RECT  159.3 309.0 160.1 308.2 ;
      RECT  162.5 309.0 163.3 308.2 ;
      RECT  160.9 309.0 161.7 308.2 ;
      RECT  160.9 315.8 161.7 315.0 ;
      RECT  159.3 315.8 160.1 315.0 ;
      RECT  162.5 315.8 163.3 315.0 ;
      RECT  160.9 315.8 161.7 315.0 ;
      RECT  159.7 312.7 160.5 311.9 ;
      RECT  161.7 314.1 162.5 313.3 ;
      RECT  163.9 312.7 164.7 311.9 ;
      RECT  158.1 307.1 165.9 306.5 ;
      RECT  158.1 317.5 165.9 316.9 ;
      RECT  168.7 309.0 169.5 308.2 ;
      RECT  167.1 309.0 167.9 308.2 ;
      RECT  168.7 316.2 169.5 315.4 ;
      RECT  167.1 316.2 167.9 315.4 ;
      RECT  167.3 312.6 168.1 311.8 ;
      RECT  169.1 312.5 169.7 311.9 ;
      RECT  165.9 307.1 172.3 306.5 ;
      RECT  165.9 317.5 172.3 316.9 ;
      RECT  167.3 312.6 168.1 311.8 ;
      RECT  169.1 312.5 169.7 311.9 ;
      RECT  165.9 307.1 166.5 306.5 ;
      RECT  165.9 317.5 166.5 316.9 ;
      RECT  160.9 325.4 161.7 326.2 ;
      RECT  159.3 325.4 160.1 326.2 ;
      RECT  162.5 325.4 163.3 326.2 ;
      RECT  160.9 325.4 161.7 326.2 ;
      RECT  160.9 318.6 161.7 319.4 ;
      RECT  159.3 318.6 160.1 319.4 ;
      RECT  162.5 318.6 163.3 319.4 ;
      RECT  160.9 318.6 161.7 319.4 ;
      RECT  159.7 321.7 160.5 322.5 ;
      RECT  161.7 320.3 162.5 321.1 ;
      RECT  163.9 321.7 164.7 322.5 ;
      RECT  158.1 327.3 165.9 327.9 ;
      RECT  158.1 316.9 165.9 317.5 ;
      RECT  168.7 325.4 169.5 326.2 ;
      RECT  167.1 325.4 167.9 326.2 ;
      RECT  168.7 318.2 169.5 319.0 ;
      RECT  167.1 318.2 167.9 319.0 ;
      RECT  167.3 321.8 168.1 322.6 ;
      RECT  169.1 321.9 169.7 322.5 ;
      RECT  165.9 327.3 172.3 327.9 ;
      RECT  165.9 316.9 172.3 317.5 ;
      RECT  167.3 321.8 168.1 322.6 ;
      RECT  169.1 321.9 169.7 322.5 ;
      RECT  165.9 327.3 166.5 327.9 ;
      RECT  165.9 316.9 166.5 317.5 ;
      RECT  160.9 329.8 161.7 329.0 ;
      RECT  159.3 329.8 160.1 329.0 ;
      RECT  162.5 329.8 163.3 329.0 ;
      RECT  160.9 329.8 161.7 329.0 ;
      RECT  160.9 336.6 161.7 335.8 ;
      RECT  159.3 336.6 160.1 335.8 ;
      RECT  162.5 336.6 163.3 335.8 ;
      RECT  160.9 336.6 161.7 335.8 ;
      RECT  159.7 333.5 160.5 332.7 ;
      RECT  161.7 334.9 162.5 334.1 ;
      RECT  163.9 333.5 164.7 332.7 ;
      RECT  158.1 327.9 165.9 327.3 ;
      RECT  158.1 338.3 165.9 337.7 ;
      RECT  168.7 329.8 169.5 329.0 ;
      RECT  167.1 329.8 167.9 329.0 ;
      RECT  168.7 337.0 169.5 336.2 ;
      RECT  167.1 337.0 167.9 336.2 ;
      RECT  167.3 333.4 168.1 332.6 ;
      RECT  169.1 333.3 169.7 332.7 ;
      RECT  165.9 327.9 172.3 327.3 ;
      RECT  165.9 338.3 172.3 337.7 ;
      RECT  167.3 333.4 168.1 332.6 ;
      RECT  169.1 333.3 169.7 332.7 ;
      RECT  165.9 327.9 166.5 327.3 ;
      RECT  165.9 338.3 166.5 337.7 ;
      RECT  160.9 346.2 161.7 347.0 ;
      RECT  159.3 346.2 160.1 347.0 ;
      RECT  162.5 346.2 163.3 347.0 ;
      RECT  160.9 346.2 161.7 347.0 ;
      RECT  160.9 339.4 161.7 340.2 ;
      RECT  159.3 339.4 160.1 340.2 ;
      RECT  162.5 339.4 163.3 340.2 ;
      RECT  160.9 339.4 161.7 340.2 ;
      RECT  159.7 342.5 160.5 343.3 ;
      RECT  161.7 341.1 162.5 341.9 ;
      RECT  163.9 342.5 164.7 343.3 ;
      RECT  158.1 348.1 165.9 348.7 ;
      RECT  158.1 337.7 165.9 338.3 ;
      RECT  168.7 346.2 169.5 347.0 ;
      RECT  167.1 346.2 167.9 347.0 ;
      RECT  168.7 339.0 169.5 339.8 ;
      RECT  167.1 339.0 167.9 339.8 ;
      RECT  167.3 342.6 168.1 343.4 ;
      RECT  169.1 342.7 169.7 343.3 ;
      RECT  165.9 348.1 172.3 348.7 ;
      RECT  165.9 337.7 172.3 338.3 ;
      RECT  167.3 342.6 168.1 343.4 ;
      RECT  169.1 342.7 169.7 343.3 ;
      RECT  165.9 348.1 166.5 348.7 ;
      RECT  165.9 337.7 166.5 338.3 ;
      RECT  160.9 350.6 161.7 349.8 ;
      RECT  159.3 350.6 160.1 349.8 ;
      RECT  162.5 350.6 163.3 349.8 ;
      RECT  160.9 350.6 161.7 349.8 ;
      RECT  160.9 357.4 161.7 356.6 ;
      RECT  159.3 357.4 160.1 356.6 ;
      RECT  162.5 357.4 163.3 356.6 ;
      RECT  160.9 357.4 161.7 356.6 ;
      RECT  159.7 354.3 160.5 353.5 ;
      RECT  161.7 355.7 162.5 354.9 ;
      RECT  163.9 354.3 164.7 353.5 ;
      RECT  158.1 348.7 165.9 348.1 ;
      RECT  158.1 359.1 165.9 358.5 ;
      RECT  168.7 350.6 169.5 349.8 ;
      RECT  167.1 350.6 167.9 349.8 ;
      RECT  168.7 357.8 169.5 357.0 ;
      RECT  167.1 357.8 167.9 357.0 ;
      RECT  167.3 354.2 168.1 353.4 ;
      RECT  169.1 354.1 169.7 353.5 ;
      RECT  165.9 348.7 172.3 348.1 ;
      RECT  165.9 359.1 172.3 358.5 ;
      RECT  167.3 354.2 168.1 353.4 ;
      RECT  169.1 354.1 169.7 353.5 ;
      RECT  165.9 348.7 166.5 348.1 ;
      RECT  165.9 359.1 166.5 358.5 ;
      RECT  153.9 195.0 157.3 195.6 ;
      RECT  153.9 210.0 157.3 210.6 ;
      RECT  153.9 215.8 157.3 216.4 ;
      RECT  153.9 230.8 157.3 231.4 ;
      RECT  153.9 236.6 157.3 237.2 ;
      RECT  153.9 251.6 157.3 252.2 ;
      RECT  153.9 257.4 157.3 258.0 ;
      RECT  153.9 272.4 157.3 273.0 ;
      RECT  153.9 278.2 157.3 278.8 ;
      RECT  153.9 293.2 157.3 293.8 ;
      RECT  153.9 299.0 157.3 299.6 ;
      RECT  153.9 314.0 157.3 314.6 ;
      RECT  153.9 319.8 157.3 320.4 ;
      RECT  153.9 334.8 157.3 335.4 ;
      RECT  153.9 340.6 157.3 341.2 ;
      RECT  153.9 355.6 157.3 356.2 ;
      RECT  169.1 197.1 169.7 197.7 ;
      RECT  169.1 207.9 169.7 208.5 ;
      RECT  169.1 217.9 169.7 218.5 ;
      RECT  169.1 228.7 169.7 229.3 ;
      RECT  169.1 238.7 169.7 239.3 ;
      RECT  169.1 249.5 169.7 250.1 ;
      RECT  169.1 259.5 169.7 260.1 ;
      RECT  169.1 270.3 169.7 270.9 ;
      RECT  169.1 280.3 169.7 280.9 ;
      RECT  169.1 291.1 169.7 291.7 ;
      RECT  169.1 301.1 169.7 301.7 ;
      RECT  169.1 311.9 169.7 312.5 ;
      RECT  169.1 321.9 169.7 322.5 ;
      RECT  169.1 332.7 169.7 333.3 ;
      RECT  169.1 342.7 169.7 343.3 ;
      RECT  169.1 353.5 169.7 354.1 ;
      RECT  169.1 197.1 169.7 197.7 ;
      RECT  169.1 207.9 169.7 208.5 ;
      RECT  169.1 217.9 169.7 218.5 ;
      RECT  169.1 228.7 169.7 229.3 ;
      RECT  169.1 238.7 169.7 239.3 ;
      RECT  169.1 249.5 169.7 250.1 ;
      RECT  169.1 259.5 169.7 260.1 ;
      RECT  169.1 270.3 169.7 270.9 ;
      RECT  169.1 280.3 169.7 280.9 ;
      RECT  169.1 291.1 169.7 291.7 ;
      RECT  169.1 301.1 169.7 301.7 ;
      RECT  169.1 311.9 169.7 312.5 ;
      RECT  169.1 321.9 169.7 322.5 ;
      RECT  169.1 332.7 169.7 333.3 ;
      RECT  169.1 342.7 169.7 343.3 ;
      RECT  169.1 353.5 169.7 354.1 ;
      RECT  1.2 10.2 11.0 10.4 ;
      RECT  15.4 9.6 19.6 10.2 ;
      RECT  18.8 1.2 19.6 5.6 ;
      RECT  7.8 13.6 11.4 14.2 ;
      RECT  18.8 6.2 19.6 9.6 ;
      RECT  7.8 4.4 8.6 4.6 ;
      RECT  10.4 12.0 12.6 12.6 ;
      RECT  1.2 1.2 2.0 6.0 ;
      RECT  11.8 6.6 12.6 6.8 ;
      RECT  7.8 13.4 8.6 13.6 ;
      RECT  4.4 12.0 5.2 12.2 ;
      RECT  11.8 11.8 12.6 12.0 ;
      RECT  12.4 10.6 14.8 11.2 ;
      RECT  5.0 7.4 5.8 7.6 ;
      RECT  18.8 10.2 19.6 18.8 ;
      RECT  15.8 5.4 16.6 5.6 ;
      RECT  14.0 8.2 17.8 8.8 ;
      RECT  6.2 4.6 6.8 6.8 ;
      RECT  8.2 0.6 9.2 3.2 ;
      RECT  17.2 0.6 18.0 5.0 ;
      RECT  9.0 12.0 9.8 12.2 ;
      RECT  17.0 8.8 17.8 9.0 ;
      RECT  10.0 14.8 10.8 18.8 ;
      RECT  4.4 14.0 5.2 14.8 ;
      RECT  14.0 14.0 14.8 14.8 ;
      RECT  6.2 10.4 11.0 10.8 ;
      RECT  1.2 10.0 7.0 10.2 ;
      RECT  3.4 8.6 8.4 9.2 ;
      RECT  10.6 13.4 11.4 13.6 ;
      RECT  4.4 14.8 6.4 15.4 ;
      RECT  2.8 0.6 3.6 5.2 ;
      RECT  7.8 3.8 10.6 4.4 ;
      RECT  20.4 0.6 21.2 2.0 ;
      RECT  1.2 10.4 2.0 18.8 ;
      RECT  2.8 11.0 3.6 19.4 ;
      RECT  14.2 11.2 14.8 12.2 ;
      RECT  14.0 2.6 15.4 3.2 ;
      RECT  8.4 14.8 9.2 19.4 ;
      RECT  11.6 14.8 12.4 19.4 ;
      RECT  14.2 12.2 15.6 13.0 ;
      RECT  12.4 7.4 13.0 10.6 ;
      RECT  2.0 6.6 3.6 6.8 ;
      RECT  4.4 2.6 6.4 3.2 ;
      RECT  5.6 1.2 6.4 2.6 ;
      RECT  14.2 14.8 15.4 18.8 ;
      RECT  6.0 3.8 6.8 4.6 ;
      RECT  10.4 10.8 11.0 12.0 ;
      RECT  7.6 9.2 8.4 9.4 ;
      RECT  14.0 8.0 14.8 8.2 ;
      RECT  10.0 14.2 10.6 14.8 ;
      RECT  4.4 11.4 9.8 12.0 ;
      RECT  10.0 1.2 10.8 3.2 ;
      RECT  0.0 19.4 21.8 20.6 ;
      RECT  5.6 15.4 6.4 18.8 ;
      RECT  17.2 10.8 18.0 19.4 ;
      RECT  1.2 9.8 6.8 10.0 ;
      RECT  3.4 8.4 4.2 8.6 ;
      RECT  11.6 0.6 12.4 3.2 ;
      RECT  14.2 1.2 15.4 2.6 ;
      RECT  0.0 -0.6 21.8 0.6 ;
      RECT  20.4 17.8 21.2 19.4 ;
      RECT  2.0 6.8 13.0 7.4 ;
      RECT  15.8 5.6 19.6 6.2 ;
      RECT  4.4 3.2 5.2 4.0 ;
      RECT  10.0 3.2 10.6 3.8 ;
      RECT  14.0 3.2 14.8 4.0 ;
      RECT  15.4 9.4 16.2 9.6 ;
      RECT  27.0 17.0 27.8 17.8 ;
      RECT  25.4 17.0 26.2 17.8 ;
      RECT  27.0 1.4 27.8 2.2 ;
      RECT  25.4 1.4 26.2 2.2 ;
      RECT  25.6 9.2 26.4 10.0 ;
      RECT  27.4 9.3 28.0 9.9 ;
      RECT  24.2 19.7 30.6 20.3 ;
      RECT  24.2 -0.3 30.6 0.3 ;
      RECT  33.4 15.4 34.2 16.2 ;
      RECT  31.8 15.4 32.6 16.2 ;
      RECT  33.4 2.2 34.2 3.0 ;
      RECT  31.8 2.2 32.6 3.0 ;
      RECT  32.0 8.8 32.8 9.6 ;
      RECT  33.8 8.9 34.4 9.5 ;
      RECT  30.6 19.7 37.0 20.3 ;
      RECT  30.6 -0.3 37.0 0.3 ;
      RECT  0.0 19.4 37.0 20.6 ;
      RECT  0.0 -0.6 37.0 0.6 ;
      RECT  1.2 29.8 11.0 29.6 ;
      RECT  15.4 30.4 19.6 29.8 ;
      RECT  18.8 38.8 19.6 34.4 ;
      RECT  7.8 26.4 11.4 25.8 ;
      RECT  18.8 33.8 19.6 30.4 ;
      RECT  7.8 35.6 8.6 35.4 ;
      RECT  10.4 28.0 12.6 27.4 ;
      RECT  1.2 38.8 2.0 34.0 ;
      RECT  11.8 33.4 12.6 33.2 ;
      RECT  7.8 26.6 8.6 26.4 ;
      RECT  4.4 28.0 5.2 27.8 ;
      RECT  11.8 28.2 12.6 28.0 ;
      RECT  12.4 29.4 14.8 28.8 ;
      RECT  5.0 32.6 5.8 32.4 ;
      RECT  18.8 29.8 19.6 21.2 ;
      RECT  15.8 34.6 16.6 34.4 ;
      RECT  14.0 31.8 17.8 31.2 ;
      RECT  6.2 35.4 6.8 33.2 ;
      RECT  8.2 39.4 9.2 36.8 ;
      RECT  17.2 39.4 18.0 35.0 ;
      RECT  9.0 28.0 9.8 27.8 ;
      RECT  17.0 31.2 17.8 31.0 ;
      RECT  10.0 25.2 10.8 21.2 ;
      RECT  4.4 26.0 5.2 25.2 ;
      RECT  14.0 26.0 14.8 25.2 ;
      RECT  6.2 29.6 11.0 29.2 ;
      RECT  1.2 30.0 7.0 29.8 ;
      RECT  3.4 31.4 8.4 30.8 ;
      RECT  10.6 26.6 11.4 26.4 ;
      RECT  4.4 25.2 6.4 24.6 ;
      RECT  2.8 39.4 3.6 34.8 ;
      RECT  7.8 36.2 10.6 35.6 ;
      RECT  20.4 39.4 21.2 38.0 ;
      RECT  1.2 29.6 2.0 21.2 ;
      RECT  2.8 29.0 3.6 20.6 ;
      RECT  14.2 28.8 14.8 27.8 ;
      RECT  14.0 37.4 15.4 36.8 ;
      RECT  8.4 25.2 9.2 20.6 ;
      RECT  11.6 25.2 12.4 20.6 ;
      RECT  14.2 27.8 15.6 27.0 ;
      RECT  12.4 32.6 13.0 29.4 ;
      RECT  2.0 33.4 3.6 33.2 ;
      RECT  4.4 37.4 6.4 36.8 ;
      RECT  5.6 38.8 6.4 37.4 ;
      RECT  14.2 25.2 15.4 21.2 ;
      RECT  6.0 36.2 6.8 35.4 ;
      RECT  10.4 29.2 11.0 28.0 ;
      RECT  7.6 30.8 8.4 30.6 ;
      RECT  14.0 32.0 14.8 31.8 ;
      RECT  10.0 25.8 10.6 25.2 ;
      RECT  4.4 28.6 9.8 28.0 ;
      RECT  10.0 38.8 10.8 36.8 ;
      RECT  0.0 20.6 21.8 19.4 ;
      RECT  5.6 24.6 6.4 21.2 ;
      RECT  17.2 29.2 18.0 20.6 ;
      RECT  1.2 30.2 6.8 30.0 ;
      RECT  3.4 31.6 4.2 31.4 ;
      RECT  11.6 39.4 12.4 36.8 ;
      RECT  14.2 38.8 15.4 37.4 ;
      RECT  0.0 40.6 21.8 39.4 ;
      RECT  20.4 22.2 21.2 20.6 ;
      RECT  2.0 33.2 13.0 32.6 ;
      RECT  15.8 34.4 19.6 33.8 ;
      RECT  4.4 36.8 5.2 36.0 ;
      RECT  10.0 36.8 10.6 36.2 ;
      RECT  14.0 36.8 14.8 36.0 ;
      RECT  15.4 30.6 16.2 30.4 ;
      RECT  27.0 23.0 27.8 22.2 ;
      RECT  25.4 23.0 26.2 22.2 ;
      RECT  27.0 38.6 27.8 37.8 ;
      RECT  25.4 38.6 26.2 37.8 ;
      RECT  25.6 30.8 26.4 30.0 ;
      RECT  27.4 30.7 28.0 30.1 ;
      RECT  24.2 20.3 30.6 19.7 ;
      RECT  24.2 40.3 30.6 39.7 ;
      RECT  33.4 24.6 34.2 23.8 ;
      RECT  31.8 24.6 32.6 23.8 ;
      RECT  33.4 37.8 34.2 37.0 ;
      RECT  31.8 37.8 32.6 37.0 ;
      RECT  32.0 31.2 32.8 30.4 ;
      RECT  33.8 31.1 34.4 30.5 ;
      RECT  30.6 20.3 37.0 19.7 ;
      RECT  30.6 40.3 37.0 39.7 ;
      RECT  0.0 20.6 37.0 19.4 ;
      RECT  0.0 40.6 37.0 39.4 ;
      RECT  52.4 17.8 53.2 18.6 ;
      RECT  50.8 17.8 51.6 18.6 ;
      RECT  52.4 1.0 53.2 1.8 ;
      RECT  50.8 1.0 51.6 1.8 ;
      RECT  51.0 9.4 51.8 10.2 ;
      RECT  52.8 9.5 53.4 10.1 ;
      RECT  49.6 19.7 56.0 20.3 ;
      RECT  49.6 -0.3 56.0 0.3 ;
      RECT  58.8 17.0 59.6 17.8 ;
      RECT  57.2 17.0 58.0 17.8 ;
      RECT  58.8 1.4 59.6 2.2 ;
      RECT  57.2 1.4 58.0 2.2 ;
      RECT  57.4 9.2 58.2 10.0 ;
      RECT  59.2 9.3 59.8 9.9 ;
      RECT  56.0 19.7 62.4 20.3 ;
      RECT  56.0 -0.3 62.4 0.3 ;
      RECT  65.2 14.6 66.0 15.4 ;
      RECT  63.6 14.6 64.4 15.4 ;
      RECT  65.2 2.6 66.0 3.4 ;
      RECT  63.6 2.6 64.4 3.4 ;
      RECT  63.8 8.6 64.6 9.4 ;
      RECT  65.6 8.7 66.2 9.3 ;
      RECT  62.4 19.7 68.8 20.3 ;
      RECT  62.4 -0.3 68.8 0.3 ;
      RECT  71.7 13.4 75.5 14.0 ;
      RECT  70.1 16.0 73.9 16.6 ;
      RECT  71.7 4.0 75.5 4.6 ;
      RECT  70.1 1.4 73.9 2.0 ;
      RECT  70.2 8.6 71.0 9.4 ;
      RECT  73.6 8.7 74.2 9.3 ;
      RECT  68.8 19.7 78.4 20.3 ;
      RECT  68.8 -0.3 78.4 0.3 ;
      RECT  51.0 9.4 51.8 10.2 ;
      RECT  73.6 8.7 74.2 9.3 ;
      RECT  49.6 19.7 50.2 20.3 ;
      RECT  49.6 -0.3 50.2 0.3 ;
      RECT  52.4 22.2 53.2 21.4 ;
      RECT  50.8 22.2 51.6 21.4 ;
      RECT  52.4 39.0 53.2 38.2 ;
      RECT  50.8 39.0 51.6 38.2 ;
      RECT  51.0 30.6 51.8 29.8 ;
      RECT  52.8 30.5 53.4 29.9 ;
      RECT  49.6 20.3 56.0 19.7 ;
      RECT  49.6 40.3 56.0 39.7 ;
      RECT  58.8 22.2 59.6 21.4 ;
      RECT  57.2 22.2 58.0 21.4 ;
      RECT  60.4 22.2 61.2 21.4 ;
      RECT  58.8 22.2 59.6 21.4 ;
      RECT  58.8 38.6 59.6 37.8 ;
      RECT  57.2 38.6 58.0 37.8 ;
      RECT  60.4 38.6 61.2 37.8 ;
      RECT  58.8 38.6 59.6 37.8 ;
      RECT  57.6 35.5 58.4 34.7 ;
      RECT  59.6 36.9 60.4 36.1 ;
      RECT  61.8 35.5 62.6 34.7 ;
      RECT  56.0 20.3 63.8 19.7 ;
      RECT  56.0 40.3 63.8 39.7 ;
      RECT  66.6 22.2 67.4 21.4 ;
      RECT  65.0 22.2 65.8 21.4 ;
      RECT  66.6 39.0 67.4 38.2 ;
      RECT  65.0 39.0 65.8 38.2 ;
      RECT  65.2 30.6 66.0 29.8 ;
      RECT  67.0 30.5 67.6 29.9 ;
      RECT  63.8 20.3 70.2 19.7 ;
      RECT  63.8 40.3 70.2 39.7 ;
      RECT  73.0 22.2 73.8 21.4 ;
      RECT  71.4 22.2 72.2 21.4 ;
      RECT  73.0 39.0 73.8 38.2 ;
      RECT  71.4 39.0 72.2 38.2 ;
      RECT  71.6 30.6 72.4 29.8 ;
      RECT  73.4 30.5 74.0 29.9 ;
      RECT  70.2 20.3 76.6 19.7 ;
      RECT  70.2 40.3 76.6 39.7 ;
      RECT  79.4 24.6 80.2 23.8 ;
      RECT  77.8 24.6 78.6 23.8 ;
      RECT  79.4 37.8 80.2 37.0 ;
      RECT  77.8 37.8 78.6 37.0 ;
      RECT  78.0 31.2 78.8 30.4 ;
      RECT  79.8 31.1 80.4 30.5 ;
      RECT  76.6 20.3 83.0 19.7 ;
      RECT  76.6 40.3 83.0 39.7 ;
      RECT  65.2 30.6 66.0 29.8 ;
      RECT  79.8 31.1 80.4 30.5 ;
      RECT  63.8 20.3 64.4 19.7 ;
      RECT  63.8 40.3 64.4 39.7 ;
      RECT  57.6 35.5 58.4 34.7 ;
      RECT  59.6 36.9 60.4 36.1 ;
      RECT  79.8 31.1 80.4 30.5 ;
      RECT  56.0 20.3 83.0 19.7 ;
      RECT  56.0 40.3 83.0 39.7 ;
      RECT  52.4 57.8 53.2 58.6 ;
      RECT  50.8 57.8 51.6 58.6 ;
      RECT  54.0 57.8 54.8 58.6 ;
      RECT  52.4 57.8 53.2 58.6 ;
      RECT  52.4 41.4 53.2 42.2 ;
      RECT  50.8 41.4 51.6 42.2 ;
      RECT  54.0 41.4 54.8 42.2 ;
      RECT  52.4 41.4 53.2 42.2 ;
      RECT  51.2 44.5 52.0 45.3 ;
      RECT  53.2 43.1 54.0 43.9 ;
      RECT  55.4 44.5 56.2 45.3 ;
      RECT  49.6 59.7 57.4 60.3 ;
      RECT  49.6 39.7 57.4 40.3 ;
      RECT  60.2 57.8 61.0 58.6 ;
      RECT  58.6 57.8 59.4 58.6 ;
      RECT  60.2 41.0 61.0 41.8 ;
      RECT  58.6 41.0 59.4 41.8 ;
      RECT  58.8 49.4 59.6 50.2 ;
      RECT  60.6 49.5 61.2 50.1 ;
      RECT  57.4 59.7 63.8 60.3 ;
      RECT  57.4 39.7 63.8 40.3 ;
      RECT  66.6 57.8 67.4 58.6 ;
      RECT  65.0 57.8 65.8 58.6 ;
      RECT  66.6 41.0 67.4 41.8 ;
      RECT  65.0 41.0 65.8 41.8 ;
      RECT  65.2 49.4 66.0 50.2 ;
      RECT  67.0 49.5 67.6 50.1 ;
      RECT  63.8 59.7 70.2 60.3 ;
      RECT  63.8 39.7 70.2 40.3 ;
      RECT  73.0 55.4 73.8 56.2 ;
      RECT  71.4 55.4 72.2 56.2 ;
      RECT  73.0 42.2 73.8 43.0 ;
      RECT  71.4 42.2 72.2 43.0 ;
      RECT  71.6 48.8 72.4 49.6 ;
      RECT  73.4 48.9 74.0 49.5 ;
      RECT  70.2 59.7 76.6 60.3 ;
      RECT  70.2 39.7 76.6 40.3 ;
      RECT  58.8 49.4 59.6 50.2 ;
      RECT  73.4 48.9 74.0 49.5 ;
      RECT  57.4 59.7 58.0 60.3 ;
      RECT  57.4 39.7 58.0 40.3 ;
      RECT  51.2 44.5 52.0 45.3 ;
      RECT  53.2 43.1 54.0 43.9 ;
      RECT  73.4 48.9 74.0 49.5 ;
      RECT  49.6 59.7 76.6 60.3 ;
      RECT  49.6 39.7 76.6 40.3 ;
      RECT  52.4 62.2 53.2 61.4 ;
      RECT  50.8 62.2 51.6 61.4 ;
      RECT  52.4 79.0 53.2 78.2 ;
      RECT  50.8 79.0 51.6 78.2 ;
      RECT  51.0 70.6 51.8 69.8 ;
      RECT  52.8 70.5 53.4 69.9 ;
      RECT  49.6 60.3 56.0 59.7 ;
      RECT  49.6 80.3 56.0 79.7 ;
      RECT  58.8 62.2 59.6 61.4 ;
      RECT  57.2 62.2 58.0 61.4 ;
      RECT  58.8 79.0 59.6 78.2 ;
      RECT  57.2 79.0 58.0 78.2 ;
      RECT  57.4 70.6 58.2 69.8 ;
      RECT  59.2 70.5 59.8 69.9 ;
      RECT  56.0 60.3 62.4 59.7 ;
      RECT  56.0 80.3 62.4 79.7 ;
      RECT  65.2 63.0 66.0 62.2 ;
      RECT  63.6 63.0 64.4 62.2 ;
      RECT  65.2 78.6 66.0 77.8 ;
      RECT  63.6 78.6 64.4 77.8 ;
      RECT  63.8 70.8 64.6 70.0 ;
      RECT  65.6 70.7 66.2 70.1 ;
      RECT  62.4 60.3 68.8 59.7 ;
      RECT  62.4 80.3 68.8 79.7 ;
      RECT  71.6 65.4 72.4 64.6 ;
      RECT  70.0 65.4 70.8 64.6 ;
      RECT  71.6 77.4 72.4 76.6 ;
      RECT  70.0 77.4 70.8 76.6 ;
      RECT  70.2 71.4 71.0 70.6 ;
      RECT  72.0 71.3 72.6 70.7 ;
      RECT  68.8 60.3 75.2 59.7 ;
      RECT  68.8 80.3 75.2 79.7 ;
      RECT  51.0 70.6 51.8 69.8 ;
      RECT  72.0 71.3 72.6 70.7 ;
      RECT  49.6 60.3 50.2 59.7 ;
      RECT  49.6 80.3 50.2 79.7 ;
      RECT  52.4 137.8 53.2 138.6 ;
      RECT  50.8 137.8 51.6 138.6 ;
      RECT  52.4 121.0 53.2 121.8 ;
      RECT  50.8 121.0 51.6 121.8 ;
      RECT  51.0 129.4 51.8 130.2 ;
      RECT  52.8 129.5 53.4 130.1 ;
      RECT  49.6 139.7 56.0 140.3 ;
      RECT  49.6 119.7 56.0 120.3 ;
      RECT  52.4 97.8 53.2 98.6 ;
      RECT  50.8 97.8 51.6 98.6 ;
      RECT  54.0 97.8 54.8 98.6 ;
      RECT  52.4 97.8 53.2 98.6 ;
      RECT  55.6 97.8 56.4 98.6 ;
      RECT  54.0 97.8 54.8 98.6 ;
      RECT  52.4 81.4 53.2 82.2 ;
      RECT  50.8 81.4 51.6 82.2 ;
      RECT  54.0 81.4 54.8 82.2 ;
      RECT  52.4 81.4 53.2 82.2 ;
      RECT  55.6 81.4 56.4 82.2 ;
      RECT  54.0 81.4 54.8 82.2 ;
      RECT  51.6 85.4 52.4 86.2 ;
      RECT  53.2 84.1 54.0 84.9 ;
      RECT  54.8 82.8 55.6 83.6 ;
      RECT  55.6 85.4 56.4 86.2 ;
      RECT  49.6 99.7 58.2 100.3 ;
      RECT  49.6 79.7 58.2 80.3 ;
      RECT  61.0 94.6 61.8 95.4 ;
      RECT  59.5 96.0 63.3 96.6 ;
      RECT  61.0 82.6 61.8 83.4 ;
      RECT  59.5 81.4 63.3 82.0 ;
      RECT  59.6 88.6 60.4 89.4 ;
      RECT  61.4 88.7 62.0 89.3 ;
      RECT  58.2 99.7 66.2 100.3 ;
      RECT  58.2 79.7 66.2 80.3 ;
      RECT  51.6 85.4 52.4 86.2 ;
      RECT  53.2 84.1 54.0 84.9 ;
      RECT  54.8 82.8 55.6 83.6 ;
      RECT  61.4 88.7 62.0 89.3 ;
      RECT  49.6 99.7 66.2 100.3 ;
      RECT  49.6 79.7 66.2 80.3 ;
      RECT  52.4 142.2 53.2 141.4 ;
      RECT  50.8 142.2 51.6 141.4 ;
      RECT  54.0 142.2 54.8 141.4 ;
      RECT  52.4 142.2 53.2 141.4 ;
      RECT  55.6 142.2 56.4 141.4 ;
      RECT  54.0 142.2 54.8 141.4 ;
      RECT  52.4 158.6 53.2 157.8 ;
      RECT  50.8 158.6 51.6 157.8 ;
      RECT  54.0 158.6 54.8 157.8 ;
      RECT  52.4 158.6 53.2 157.8 ;
      RECT  55.6 158.6 56.4 157.8 ;
      RECT  54.0 158.6 54.8 157.8 ;
      RECT  51.6 154.6 52.4 153.8 ;
      RECT  53.2 155.9 54.0 155.1 ;
      RECT  54.8 157.2 55.6 156.4 ;
      RECT  55.6 154.6 56.4 153.8 ;
      RECT  49.6 140.3 58.2 139.7 ;
      RECT  49.6 160.3 58.2 159.7 ;
      RECT  61.0 143.0 61.8 142.2 ;
      RECT  59.4 143.0 60.2 142.2 ;
      RECT  61.0 158.6 61.8 157.8 ;
      RECT  59.4 158.6 60.2 157.8 ;
      RECT  59.6 150.8 60.4 150.0 ;
      RECT  61.4 150.7 62.0 150.1 ;
      RECT  58.2 140.3 64.6 139.7 ;
      RECT  58.2 160.3 64.6 159.7 ;
      RECT  51.6 154.6 52.4 153.8 ;
      RECT  53.2 155.9 54.0 155.1 ;
      RECT  54.8 157.2 55.6 156.4 ;
      RECT  61.4 150.7 62.0 150.1 ;
      RECT  49.6 140.3 64.6 139.7 ;
      RECT  49.6 160.3 64.6 159.7 ;
      RECT  29.2 171.8 28.4 172.6 ;
      RECT  30.8 171.8 30.0 172.6 ;
      RECT  29.2 163.8 28.4 164.6 ;
      RECT  30.8 163.8 30.0 164.6 ;
      RECT  30.6 167.8 29.8 168.6 ;
      RECT  28.8 167.9 28.2 168.5 ;
      RECT  32.0 173.7 25.6 174.3 ;
      RECT  32.0 162.5 25.6 163.1 ;
      RECT  22.8 171.8 22.0 172.6 ;
      RECT  24.4 171.8 23.6 172.6 ;
      RECT  22.8 163.8 22.0 164.6 ;
      RECT  24.4 163.8 23.6 164.6 ;
      RECT  24.2 167.8 23.4 168.6 ;
      RECT  22.4 167.9 21.8 168.5 ;
      RECT  25.6 173.7 19.2 174.3 ;
      RECT  25.6 162.5 19.2 163.1 ;
      RECT  16.4 171.8 15.6 172.6 ;
      RECT  18.0 171.8 17.2 172.6 ;
      RECT  16.4 163.8 15.6 164.6 ;
      RECT  18.0 163.8 17.2 164.6 ;
      RECT  17.8 167.8 17.0 168.6 ;
      RECT  16.0 167.9 15.4 168.5 ;
      RECT  19.2 173.7 12.8 174.3 ;
      RECT  19.2 162.5 12.8 163.1 ;
      RECT  10.0 171.8 9.2 172.6 ;
      RECT  11.6 171.8 10.8 172.6 ;
      RECT  10.0 163.8 9.2 164.6 ;
      RECT  11.6 163.8 10.8 164.6 ;
      RECT  11.4 167.8 10.6 168.6 ;
      RECT  9.6 167.9 9.0 168.5 ;
      RECT  12.8 173.7 6.4 174.3 ;
      RECT  12.8 162.5 6.4 163.1 ;
      RECT  3.6 171.8 2.8 172.6 ;
      RECT  5.2 171.8 4.4 172.6 ;
      RECT  3.6 163.8 2.8 164.6 ;
      RECT  5.2 163.8 4.4 164.6 ;
      RECT  5.0 167.8 4.2 168.6 ;
      RECT  3.2 167.9 2.6 168.5 ;
      RECT  6.4 173.7 0.0 174.3 ;
      RECT  6.4 162.5 0.0 163.1 ;
      RECT  29.2 176.2 28.4 175.4 ;
      RECT  30.8 176.2 30.0 175.4 ;
      RECT  29.2 184.2 28.4 183.4 ;
      RECT  30.8 184.2 30.0 183.4 ;
      RECT  30.6 180.2 29.8 179.4 ;
      RECT  28.8 180.1 28.2 179.5 ;
      RECT  32.0 174.3 25.6 173.7 ;
      RECT  32.0 185.5 25.6 184.9 ;
      RECT  22.8 176.2 22.0 175.4 ;
      RECT  24.4 176.2 23.6 175.4 ;
      RECT  22.8 184.2 22.0 183.4 ;
      RECT  24.4 184.2 23.6 183.4 ;
      RECT  24.2 180.2 23.4 179.4 ;
      RECT  22.4 180.1 21.8 179.5 ;
      RECT  25.6 174.3 19.2 173.7 ;
      RECT  25.6 185.5 19.2 184.9 ;
      RECT  16.4 176.2 15.6 175.4 ;
      RECT  18.0 176.2 17.2 175.4 ;
      RECT  16.4 184.2 15.6 183.4 ;
      RECT  18.0 184.2 17.2 183.4 ;
      RECT  17.8 180.2 17.0 179.4 ;
      RECT  16.0 180.1 15.4 179.5 ;
      RECT  19.2 174.3 12.8 173.7 ;
      RECT  19.2 185.5 12.8 184.9 ;
      RECT  10.0 176.2 9.2 175.4 ;
      RECT  11.6 176.2 10.8 175.4 ;
      RECT  10.0 184.2 9.2 183.4 ;
      RECT  11.6 184.2 10.8 183.4 ;
      RECT  11.4 180.2 10.6 179.4 ;
      RECT  9.6 180.1 9.0 179.5 ;
      RECT  12.8 174.3 6.4 173.7 ;
      RECT  12.8 185.5 6.4 184.9 ;
      RECT  3.6 176.2 2.8 175.4 ;
      RECT  5.2 176.2 4.4 175.4 ;
      RECT  3.6 184.2 2.8 183.4 ;
      RECT  5.2 184.2 4.4 183.4 ;
      RECT  5.0 180.2 4.2 179.4 ;
      RECT  3.2 180.1 2.6 179.5 ;
      RECT  6.4 174.3 0.0 173.7 ;
      RECT  6.4 185.5 0.0 184.9 ;
      RECT  29.2 194.2 28.4 195.0 ;
      RECT  30.8 194.2 30.0 195.0 ;
      RECT  29.2 186.2 28.4 187.0 ;
      RECT  30.8 186.2 30.0 187.0 ;
      RECT  30.6 190.2 29.8 191.0 ;
      RECT  28.8 190.3 28.2 190.9 ;
      RECT  32.0 196.1 25.6 196.7 ;
      RECT  32.0 184.9 25.6 185.5 ;
      RECT  22.8 194.2 22.0 195.0 ;
      RECT  24.4 194.2 23.6 195.0 ;
      RECT  22.8 186.2 22.0 187.0 ;
      RECT  24.4 186.2 23.6 187.0 ;
      RECT  24.2 190.2 23.4 191.0 ;
      RECT  22.4 190.3 21.8 190.9 ;
      RECT  25.6 196.1 19.2 196.7 ;
      RECT  25.6 184.9 19.2 185.5 ;
      RECT  16.4 194.2 15.6 195.0 ;
      RECT  18.0 194.2 17.2 195.0 ;
      RECT  16.4 186.2 15.6 187.0 ;
      RECT  18.0 186.2 17.2 187.0 ;
      RECT  17.8 190.2 17.0 191.0 ;
      RECT  16.0 190.3 15.4 190.9 ;
      RECT  19.2 196.1 12.8 196.7 ;
      RECT  19.2 184.9 12.8 185.5 ;
      RECT  10.0 194.2 9.2 195.0 ;
      RECT  11.6 194.2 10.8 195.0 ;
      RECT  10.0 186.2 9.2 187.0 ;
      RECT  11.6 186.2 10.8 187.0 ;
      RECT  11.4 190.2 10.6 191.0 ;
      RECT  9.6 190.3 9.0 190.9 ;
      RECT  12.8 196.1 6.4 196.7 ;
      RECT  12.8 184.9 6.4 185.5 ;
      RECT  3.6 194.2 2.8 195.0 ;
      RECT  5.2 194.2 4.4 195.0 ;
      RECT  3.6 186.2 2.8 187.0 ;
      RECT  5.2 186.2 4.4 187.0 ;
      RECT  5.0 190.2 4.2 191.0 ;
      RECT  3.2 190.3 2.6 190.9 ;
      RECT  6.4 196.1 0.0 196.7 ;
      RECT  6.4 184.9 0.0 185.5 ;
      RECT  29.2 198.6 28.4 197.8 ;
      RECT  30.8 198.6 30.0 197.8 ;
      RECT  29.2 206.6 28.4 205.8 ;
      RECT  30.8 206.6 30.0 205.8 ;
      RECT  30.6 202.6 29.8 201.8 ;
      RECT  28.8 202.5 28.2 201.9 ;
      RECT  32.0 196.7 25.6 196.1 ;
      RECT  32.0 207.9 25.6 207.3 ;
      RECT  22.8 198.6 22.0 197.8 ;
      RECT  24.4 198.6 23.6 197.8 ;
      RECT  22.8 206.6 22.0 205.8 ;
      RECT  24.4 206.6 23.6 205.8 ;
      RECT  24.2 202.6 23.4 201.8 ;
      RECT  22.4 202.5 21.8 201.9 ;
      RECT  25.6 196.7 19.2 196.1 ;
      RECT  25.6 207.9 19.2 207.3 ;
      RECT  16.4 198.6 15.6 197.8 ;
      RECT  18.0 198.6 17.2 197.8 ;
      RECT  16.4 206.6 15.6 205.8 ;
      RECT  18.0 206.6 17.2 205.8 ;
      RECT  17.8 202.6 17.0 201.8 ;
      RECT  16.0 202.5 15.4 201.9 ;
      RECT  19.2 196.7 12.8 196.1 ;
      RECT  19.2 207.9 12.8 207.3 ;
      RECT  10.0 198.6 9.2 197.8 ;
      RECT  11.6 198.6 10.8 197.8 ;
      RECT  10.0 206.6 9.2 205.8 ;
      RECT  11.6 206.6 10.8 205.8 ;
      RECT  11.4 202.6 10.6 201.8 ;
      RECT  9.6 202.5 9.0 201.9 ;
      RECT  12.8 196.7 6.4 196.1 ;
      RECT  12.8 207.9 6.4 207.3 ;
      RECT  3.6 198.6 2.8 197.8 ;
      RECT  5.2 198.6 4.4 197.8 ;
      RECT  3.6 206.6 2.8 205.8 ;
      RECT  5.2 206.6 4.4 205.8 ;
      RECT  5.0 202.6 4.2 201.8 ;
      RECT  3.2 202.5 2.6 201.9 ;
      RECT  6.4 196.7 0.0 196.1 ;
      RECT  6.4 207.9 0.0 207.3 ;
      RECT  29.2 216.6 28.4 217.4 ;
      RECT  30.8 216.6 30.0 217.4 ;
      RECT  29.2 208.6 28.4 209.4 ;
      RECT  30.8 208.6 30.0 209.4 ;
      RECT  30.6 212.6 29.8 213.4 ;
      RECT  28.8 212.7 28.2 213.3 ;
      RECT  32.0 218.5 25.6 219.1 ;
      RECT  32.0 207.3 25.6 207.9 ;
      RECT  22.8 216.6 22.0 217.4 ;
      RECT  24.4 216.6 23.6 217.4 ;
      RECT  22.8 208.6 22.0 209.4 ;
      RECT  24.4 208.6 23.6 209.4 ;
      RECT  24.2 212.6 23.4 213.4 ;
      RECT  22.4 212.7 21.8 213.3 ;
      RECT  25.6 218.5 19.2 219.1 ;
      RECT  25.6 207.3 19.2 207.9 ;
      RECT  16.4 216.6 15.6 217.4 ;
      RECT  18.0 216.6 17.2 217.4 ;
      RECT  16.4 208.6 15.6 209.4 ;
      RECT  18.0 208.6 17.2 209.4 ;
      RECT  17.8 212.6 17.0 213.4 ;
      RECT  16.0 212.7 15.4 213.3 ;
      RECT  19.2 218.5 12.8 219.1 ;
      RECT  19.2 207.3 12.8 207.9 ;
      RECT  10.0 216.6 9.2 217.4 ;
      RECT  11.6 216.6 10.8 217.4 ;
      RECT  10.0 208.6 9.2 209.4 ;
      RECT  11.6 208.6 10.8 209.4 ;
      RECT  11.4 212.6 10.6 213.4 ;
      RECT  9.6 212.7 9.0 213.3 ;
      RECT  12.8 218.5 6.4 219.1 ;
      RECT  12.8 207.3 6.4 207.9 ;
      RECT  3.6 216.6 2.8 217.4 ;
      RECT  5.2 216.6 4.4 217.4 ;
      RECT  3.6 208.6 2.8 209.4 ;
      RECT  5.2 208.6 4.4 209.4 ;
      RECT  5.0 212.6 4.2 213.4 ;
      RECT  3.2 212.7 2.6 213.3 ;
      RECT  6.4 218.5 0.0 219.1 ;
      RECT  6.4 207.3 0.0 207.9 ;
      RECT  29.2 221.0 28.4 220.2 ;
      RECT  30.8 221.0 30.0 220.2 ;
      RECT  29.2 229.0 28.4 228.2 ;
      RECT  30.8 229.0 30.0 228.2 ;
      RECT  30.6 225.0 29.8 224.2 ;
      RECT  28.8 224.9 28.2 224.3 ;
      RECT  32.0 219.1 25.6 218.5 ;
      RECT  32.0 230.3 25.6 229.7 ;
      RECT  22.8 221.0 22.0 220.2 ;
      RECT  24.4 221.0 23.6 220.2 ;
      RECT  22.8 229.0 22.0 228.2 ;
      RECT  24.4 229.0 23.6 228.2 ;
      RECT  24.2 225.0 23.4 224.2 ;
      RECT  22.4 224.9 21.8 224.3 ;
      RECT  25.6 219.1 19.2 218.5 ;
      RECT  25.6 230.3 19.2 229.7 ;
      RECT  16.4 221.0 15.6 220.2 ;
      RECT  18.0 221.0 17.2 220.2 ;
      RECT  16.4 229.0 15.6 228.2 ;
      RECT  18.0 229.0 17.2 228.2 ;
      RECT  17.8 225.0 17.0 224.2 ;
      RECT  16.0 224.9 15.4 224.3 ;
      RECT  19.2 219.1 12.8 218.5 ;
      RECT  19.2 230.3 12.8 229.7 ;
      RECT  10.0 221.0 9.2 220.2 ;
      RECT  11.6 221.0 10.8 220.2 ;
      RECT  10.0 229.0 9.2 228.2 ;
      RECT  11.6 229.0 10.8 228.2 ;
      RECT  11.4 225.0 10.6 224.2 ;
      RECT  9.6 224.9 9.0 224.3 ;
      RECT  12.8 219.1 6.4 218.5 ;
      RECT  12.8 230.3 6.4 229.7 ;
      RECT  3.6 221.0 2.8 220.2 ;
      RECT  5.2 221.0 4.4 220.2 ;
      RECT  3.6 229.0 2.8 228.2 ;
      RECT  5.2 229.0 4.4 228.2 ;
      RECT  5.0 225.0 4.2 224.2 ;
      RECT  3.2 224.9 2.6 224.3 ;
      RECT  6.4 219.1 0.0 218.5 ;
      RECT  6.4 230.3 0.0 229.7 ;
      RECT  29.2 239.0 28.4 239.8 ;
      RECT  30.8 239.0 30.0 239.8 ;
      RECT  29.2 231.0 28.4 231.8 ;
      RECT  30.8 231.0 30.0 231.8 ;
      RECT  30.6 235.0 29.8 235.8 ;
      RECT  28.8 235.1 28.2 235.7 ;
      RECT  32.0 240.9 25.6 241.5 ;
      RECT  32.0 229.7 25.6 230.3 ;
      RECT  22.8 239.0 22.0 239.8 ;
      RECT  24.4 239.0 23.6 239.8 ;
      RECT  22.8 231.0 22.0 231.8 ;
      RECT  24.4 231.0 23.6 231.8 ;
      RECT  24.2 235.0 23.4 235.8 ;
      RECT  22.4 235.1 21.8 235.7 ;
      RECT  25.6 240.9 19.2 241.5 ;
      RECT  25.6 229.7 19.2 230.3 ;
      RECT  16.4 239.0 15.6 239.8 ;
      RECT  18.0 239.0 17.2 239.8 ;
      RECT  16.4 231.0 15.6 231.8 ;
      RECT  18.0 231.0 17.2 231.8 ;
      RECT  17.8 235.0 17.0 235.8 ;
      RECT  16.0 235.1 15.4 235.7 ;
      RECT  19.2 240.9 12.8 241.5 ;
      RECT  19.2 229.7 12.8 230.3 ;
      RECT  10.0 239.0 9.2 239.8 ;
      RECT  11.6 239.0 10.8 239.8 ;
      RECT  10.0 231.0 9.2 231.8 ;
      RECT  11.6 231.0 10.8 231.8 ;
      RECT  11.4 235.0 10.6 235.8 ;
      RECT  9.6 235.1 9.0 235.7 ;
      RECT  12.8 240.9 6.4 241.5 ;
      RECT  12.8 229.7 6.4 230.3 ;
      RECT  3.6 239.0 2.8 239.8 ;
      RECT  5.2 239.0 4.4 239.8 ;
      RECT  3.6 231.0 2.8 231.8 ;
      RECT  5.2 231.0 4.4 231.8 ;
      RECT  5.0 235.0 4.2 235.8 ;
      RECT  3.2 235.1 2.6 235.7 ;
      RECT  6.4 240.9 0.0 241.5 ;
      RECT  6.4 229.7 0.0 230.3 ;
      RECT  29.2 243.4 28.4 242.6 ;
      RECT  30.8 243.4 30.0 242.6 ;
      RECT  29.2 251.4 28.4 250.6 ;
      RECT  30.8 251.4 30.0 250.6 ;
      RECT  30.6 247.4 29.8 246.6 ;
      RECT  28.8 247.3 28.2 246.7 ;
      RECT  32.0 241.5 25.6 240.9 ;
      RECT  32.0 252.7 25.6 252.1 ;
      RECT  22.8 243.4 22.0 242.6 ;
      RECT  24.4 243.4 23.6 242.6 ;
      RECT  22.8 251.4 22.0 250.6 ;
      RECT  24.4 251.4 23.6 250.6 ;
      RECT  24.2 247.4 23.4 246.6 ;
      RECT  22.4 247.3 21.8 246.7 ;
      RECT  25.6 241.5 19.2 240.9 ;
      RECT  25.6 252.7 19.2 252.1 ;
      RECT  16.4 243.4 15.6 242.6 ;
      RECT  18.0 243.4 17.2 242.6 ;
      RECT  16.4 251.4 15.6 250.6 ;
      RECT  18.0 251.4 17.2 250.6 ;
      RECT  17.8 247.4 17.0 246.6 ;
      RECT  16.0 247.3 15.4 246.7 ;
      RECT  19.2 241.5 12.8 240.9 ;
      RECT  19.2 252.7 12.8 252.1 ;
      RECT  10.0 243.4 9.2 242.6 ;
      RECT  11.6 243.4 10.8 242.6 ;
      RECT  10.0 251.4 9.2 250.6 ;
      RECT  11.6 251.4 10.8 250.6 ;
      RECT  11.4 247.4 10.6 246.6 ;
      RECT  9.6 247.3 9.0 246.7 ;
      RECT  12.8 241.5 6.4 240.9 ;
      RECT  12.8 252.7 6.4 252.1 ;
      RECT  3.6 243.4 2.8 242.6 ;
      RECT  5.2 243.4 4.4 242.6 ;
      RECT  3.6 251.4 2.8 250.6 ;
      RECT  5.2 251.4 4.4 250.6 ;
      RECT  5.0 247.4 4.2 246.6 ;
      RECT  3.2 247.3 2.6 246.7 ;
      RECT  6.4 241.5 0.0 240.9 ;
      RECT  6.4 252.7 0.0 252.1 ;
      RECT  29.2 261.4 28.4 262.2 ;
      RECT  30.8 261.4 30.0 262.2 ;
      RECT  29.2 253.4 28.4 254.2 ;
      RECT  30.8 253.4 30.0 254.2 ;
      RECT  30.6 257.4 29.8 258.2 ;
      RECT  28.8 257.5 28.2 258.1 ;
      RECT  32.0 263.3 25.6 263.9 ;
      RECT  32.0 252.1 25.6 252.7 ;
      RECT  22.8 261.4 22.0 262.2 ;
      RECT  24.4 261.4 23.6 262.2 ;
      RECT  22.8 253.4 22.0 254.2 ;
      RECT  24.4 253.4 23.6 254.2 ;
      RECT  24.2 257.4 23.4 258.2 ;
      RECT  22.4 257.5 21.8 258.1 ;
      RECT  25.6 263.3 19.2 263.9 ;
      RECT  25.6 252.1 19.2 252.7 ;
      RECT  16.4 261.4 15.6 262.2 ;
      RECT  18.0 261.4 17.2 262.2 ;
      RECT  16.4 253.4 15.6 254.2 ;
      RECT  18.0 253.4 17.2 254.2 ;
      RECT  17.8 257.4 17.0 258.2 ;
      RECT  16.0 257.5 15.4 258.1 ;
      RECT  19.2 263.3 12.8 263.9 ;
      RECT  19.2 252.1 12.8 252.7 ;
      RECT  10.0 261.4 9.2 262.2 ;
      RECT  11.6 261.4 10.8 262.2 ;
      RECT  10.0 253.4 9.2 254.2 ;
      RECT  11.6 253.4 10.8 254.2 ;
      RECT  11.4 257.4 10.6 258.2 ;
      RECT  9.6 257.5 9.0 258.1 ;
      RECT  12.8 263.3 6.4 263.9 ;
      RECT  12.8 252.1 6.4 252.7 ;
      RECT  3.6 261.4 2.8 262.2 ;
      RECT  5.2 261.4 4.4 262.2 ;
      RECT  3.6 253.4 2.8 254.2 ;
      RECT  5.2 253.4 4.4 254.2 ;
      RECT  5.0 257.4 4.2 258.2 ;
      RECT  3.2 257.5 2.6 258.1 ;
      RECT  6.4 263.3 0.0 263.9 ;
      RECT  6.4 252.1 0.0 252.7 ;
      RECT  52.4 102.2 53.2 101.4 ;
      RECT  50.8 102.2 51.6 101.4 ;
      RECT  54.0 102.2 54.8 101.4 ;
      RECT  52.4 102.2 53.2 101.4 ;
      RECT  52.4 118.6 53.2 117.8 ;
      RECT  50.8 118.6 51.6 117.8 ;
      RECT  54.0 118.6 54.8 117.8 ;
      RECT  52.4 118.6 53.2 117.8 ;
      RECT  51.2 115.5 52.0 114.7 ;
      RECT  53.2 116.9 54.0 116.1 ;
      RECT  55.4 115.5 56.2 114.7 ;
      RECT  49.6 100.3 57.4 99.7 ;
      RECT  49.6 120.3 57.4 119.7 ;
      RECT  60.2 102.2 61.0 101.4 ;
      RECT  58.6 102.2 59.4 101.4 ;
      RECT  60.2 119.0 61.0 118.2 ;
      RECT  58.6 119.0 59.4 118.2 ;
      RECT  58.8 110.6 59.6 109.8 ;
      RECT  60.6 110.5 61.2 109.9 ;
      RECT  57.4 100.3 63.8 99.7 ;
      RECT  57.4 120.3 63.8 119.7 ;
      RECT  66.6 102.2 67.4 101.4 ;
      RECT  65.0 102.2 65.8 101.4 ;
      RECT  66.6 119.0 67.4 118.2 ;
      RECT  65.0 119.0 65.8 118.2 ;
      RECT  65.2 110.6 66.0 109.8 ;
      RECT  67.0 110.5 67.6 109.9 ;
      RECT  63.8 100.3 70.2 99.7 ;
      RECT  63.8 120.3 70.2 119.7 ;
      RECT  58.8 110.6 59.6 109.8 ;
      RECT  67.0 110.5 67.6 109.9 ;
      RECT  57.4 100.3 58.0 99.7 ;
      RECT  57.4 120.3 58.0 119.7 ;
      RECT  61.7 150.1 84.4 150.7 ;
      RECT  61.7 88.7 84.4 89.3 ;
      RECT  67.3 109.9 84.4 110.5 ;
      RECT  72.3 70.7 84.4 71.3 ;
      RECT  73.9 8.7 84.4 9.3 ;
      RECT  63.8 300.8 73.6 301.0 ;
      RECT  78.0 300.2 82.2 300.8 ;
      RECT  81.4 291.8 82.2 296.2 ;
      RECT  70.4 304.2 74.0 304.8 ;
      RECT  81.4 296.8 82.2 300.2 ;
      RECT  70.4 295.0 71.2 295.2 ;
      RECT  73.0 302.6 75.2 303.2 ;
      RECT  63.8 291.8 64.6 296.6 ;
      RECT  74.4 297.2 75.2 297.4 ;
      RECT  70.4 304.0 71.2 304.2 ;
      RECT  67.0 302.6 67.8 302.8 ;
      RECT  74.4 302.4 75.2 302.6 ;
      RECT  75.0 301.2 77.4 301.8 ;
      RECT  67.6 298.0 68.4 298.2 ;
      RECT  81.4 300.8 82.2 309.4 ;
      RECT  78.4 296.0 79.2 296.2 ;
      RECT  76.6 298.8 80.4 299.4 ;
      RECT  68.8 295.2 69.4 297.4 ;
      RECT  70.8 291.2 71.8 293.8 ;
      RECT  79.8 291.2 80.6 295.6 ;
      RECT  71.6 302.6 72.4 302.8 ;
      RECT  79.6 299.4 80.4 299.6 ;
      RECT  72.6 305.4 73.4 309.4 ;
      RECT  67.0 304.6 67.8 305.4 ;
      RECT  76.6 304.6 77.4 305.4 ;
      RECT  68.8 301.0 73.6 301.4 ;
      RECT  63.8 300.6 69.6 300.8 ;
      RECT  66.0 299.2 71.0 299.8 ;
      RECT  73.2 304.0 74.0 304.2 ;
      RECT  67.0 305.4 69.0 306.0 ;
      RECT  65.4 291.2 66.2 295.8 ;
      RECT  70.4 294.4 73.2 295.0 ;
      RECT  83.0 291.2 83.8 292.6 ;
      RECT  63.8 301.0 64.6 309.4 ;
      RECT  65.4 301.6 66.2 310.0 ;
      RECT  76.8 301.8 77.4 302.8 ;
      RECT  76.6 293.2 78.0 293.8 ;
      RECT  71.0 305.4 71.8 310.0 ;
      RECT  74.2 305.4 75.0 310.0 ;
      RECT  76.8 302.8 78.2 303.6 ;
      RECT  75.0 298.0 75.6 301.2 ;
      RECT  64.6 297.2 66.2 297.4 ;
      RECT  67.0 293.2 69.0 293.8 ;
      RECT  68.2 291.8 69.0 293.2 ;
      RECT  76.8 305.4 78.0 309.4 ;
      RECT  68.6 294.4 69.4 295.2 ;
      RECT  73.0 301.4 73.6 302.6 ;
      RECT  70.2 299.8 71.0 300.0 ;
      RECT  76.6 298.6 77.4 298.8 ;
      RECT  72.6 304.8 73.2 305.4 ;
      RECT  67.0 302.0 72.4 302.6 ;
      RECT  72.6 291.8 73.4 293.8 ;
      RECT  62.6 310.0 84.4 311.2 ;
      RECT  68.2 306.0 69.0 309.4 ;
      RECT  79.8 301.4 80.6 310.0 ;
      RECT  63.8 300.4 69.4 300.6 ;
      RECT  66.0 299.0 66.8 299.2 ;
      RECT  74.2 291.2 75.0 293.8 ;
      RECT  76.8 291.8 78.0 293.2 ;
      RECT  62.6 290.0 84.4 291.2 ;
      RECT  83.0 308.4 83.8 310.0 ;
      RECT  64.6 297.4 75.6 298.0 ;
      RECT  78.4 296.2 82.2 296.8 ;
      RECT  67.0 293.8 67.8 294.6 ;
      RECT  72.6 293.8 73.2 294.4 ;
      RECT  76.6 293.8 77.4 294.6 ;
      RECT  78.0 300.0 78.8 300.2 ;
      RECT  63.8 320.4 73.6 320.2 ;
      RECT  78.0 321.0 82.2 320.4 ;
      RECT  81.4 329.4 82.2 325.0 ;
      RECT  70.4 317.0 74.0 316.4 ;
      RECT  81.4 324.4 82.2 321.0 ;
      RECT  70.4 326.2 71.2 326.0 ;
      RECT  73.0 318.6 75.2 318.0 ;
      RECT  63.8 329.4 64.6 324.6 ;
      RECT  74.4 324.0 75.2 323.8 ;
      RECT  70.4 317.2 71.2 317.0 ;
      RECT  67.0 318.6 67.8 318.4 ;
      RECT  74.4 318.8 75.2 318.6 ;
      RECT  75.0 320.0 77.4 319.4 ;
      RECT  67.6 323.2 68.4 323.0 ;
      RECT  81.4 320.4 82.2 311.8 ;
      RECT  78.4 325.2 79.2 325.0 ;
      RECT  76.6 322.4 80.4 321.8 ;
      RECT  68.8 326.0 69.4 323.8 ;
      RECT  70.8 330.0 71.8 327.4 ;
      RECT  79.8 330.0 80.6 325.6 ;
      RECT  71.6 318.6 72.4 318.4 ;
      RECT  79.6 321.8 80.4 321.6 ;
      RECT  72.6 315.8 73.4 311.8 ;
      RECT  67.0 316.6 67.8 315.8 ;
      RECT  76.6 316.6 77.4 315.8 ;
      RECT  68.8 320.2 73.6 319.8 ;
      RECT  63.8 320.6 69.6 320.4 ;
      RECT  66.0 322.0 71.0 321.4 ;
      RECT  73.2 317.2 74.0 317.0 ;
      RECT  67.0 315.8 69.0 315.2 ;
      RECT  65.4 330.0 66.2 325.4 ;
      RECT  70.4 326.8 73.2 326.2 ;
      RECT  83.0 330.0 83.8 328.6 ;
      RECT  63.8 320.2 64.6 311.8 ;
      RECT  65.4 319.6 66.2 311.2 ;
      RECT  76.8 319.4 77.4 318.4 ;
      RECT  76.6 328.0 78.0 327.4 ;
      RECT  71.0 315.8 71.8 311.2 ;
      RECT  74.2 315.8 75.0 311.2 ;
      RECT  76.8 318.4 78.2 317.6 ;
      RECT  75.0 323.2 75.6 320.0 ;
      RECT  64.6 324.0 66.2 323.8 ;
      RECT  67.0 328.0 69.0 327.4 ;
      RECT  68.2 329.4 69.0 328.0 ;
      RECT  76.8 315.8 78.0 311.8 ;
      RECT  68.6 326.8 69.4 326.0 ;
      RECT  73.0 319.8 73.6 318.6 ;
      RECT  70.2 321.4 71.0 321.2 ;
      RECT  76.6 322.6 77.4 322.4 ;
      RECT  72.6 316.4 73.2 315.8 ;
      RECT  67.0 319.2 72.4 318.6 ;
      RECT  72.6 329.4 73.4 327.4 ;
      RECT  62.6 311.2 84.4 310.0 ;
      RECT  68.2 315.2 69.0 311.8 ;
      RECT  79.8 319.8 80.6 311.2 ;
      RECT  63.8 320.8 69.4 320.6 ;
      RECT  66.0 322.2 66.8 322.0 ;
      RECT  74.2 330.0 75.0 327.4 ;
      RECT  76.8 329.4 78.0 328.0 ;
      RECT  62.6 331.2 84.4 330.0 ;
      RECT  83.0 312.8 83.8 311.2 ;
      RECT  64.6 323.8 75.6 323.2 ;
      RECT  78.4 325.0 82.2 324.4 ;
      RECT  67.0 327.4 67.8 326.6 ;
      RECT  72.6 327.4 73.2 326.8 ;
      RECT  76.6 327.4 77.4 326.6 ;
      RECT  78.0 321.2 78.8 321.0 ;
      RECT  63.8 340.8 73.6 341.0 ;
      RECT  78.0 340.2 82.2 340.8 ;
      RECT  81.4 331.8 82.2 336.2 ;
      RECT  70.4 344.2 74.0 344.8 ;
      RECT  81.4 336.8 82.2 340.2 ;
      RECT  70.4 335.0 71.2 335.2 ;
      RECT  73.0 342.6 75.2 343.2 ;
      RECT  63.8 331.8 64.6 336.6 ;
      RECT  74.4 337.2 75.2 337.4 ;
      RECT  70.4 344.0 71.2 344.2 ;
      RECT  67.0 342.6 67.8 342.8 ;
      RECT  74.4 342.4 75.2 342.6 ;
      RECT  75.0 341.2 77.4 341.8 ;
      RECT  67.6 338.0 68.4 338.2 ;
      RECT  81.4 340.8 82.2 349.4 ;
      RECT  78.4 336.0 79.2 336.2 ;
      RECT  76.6 338.8 80.4 339.4 ;
      RECT  68.8 335.2 69.4 337.4 ;
      RECT  70.8 331.2 71.8 333.8 ;
      RECT  79.8 331.2 80.6 335.6 ;
      RECT  71.6 342.6 72.4 342.8 ;
      RECT  79.6 339.4 80.4 339.6 ;
      RECT  72.6 345.4 73.4 349.4 ;
      RECT  67.0 344.6 67.8 345.4 ;
      RECT  76.6 344.6 77.4 345.4 ;
      RECT  68.8 341.0 73.6 341.4 ;
      RECT  63.8 340.6 69.6 340.8 ;
      RECT  66.0 339.2 71.0 339.8 ;
      RECT  73.2 344.0 74.0 344.2 ;
      RECT  67.0 345.4 69.0 346.0 ;
      RECT  65.4 331.2 66.2 335.8 ;
      RECT  70.4 334.4 73.2 335.0 ;
      RECT  83.0 331.2 83.8 332.6 ;
      RECT  63.8 341.0 64.6 349.4 ;
      RECT  65.4 341.6 66.2 350.0 ;
      RECT  76.8 341.8 77.4 342.8 ;
      RECT  76.6 333.2 78.0 333.8 ;
      RECT  71.0 345.4 71.8 350.0 ;
      RECT  74.2 345.4 75.0 350.0 ;
      RECT  76.8 342.8 78.2 343.6 ;
      RECT  75.0 338.0 75.6 341.2 ;
      RECT  64.6 337.2 66.2 337.4 ;
      RECT  67.0 333.2 69.0 333.8 ;
      RECT  68.2 331.8 69.0 333.2 ;
      RECT  76.8 345.4 78.0 349.4 ;
      RECT  68.6 334.4 69.4 335.2 ;
      RECT  73.0 341.4 73.6 342.6 ;
      RECT  70.2 339.8 71.0 340.0 ;
      RECT  76.6 338.6 77.4 338.8 ;
      RECT  72.6 344.8 73.2 345.4 ;
      RECT  67.0 342.0 72.4 342.6 ;
      RECT  72.6 331.8 73.4 333.8 ;
      RECT  62.6 350.0 84.4 351.2 ;
      RECT  68.2 346.0 69.0 349.4 ;
      RECT  79.8 341.4 80.6 350.0 ;
      RECT  63.8 340.4 69.4 340.6 ;
      RECT  66.0 339.0 66.8 339.2 ;
      RECT  74.2 331.2 75.0 333.8 ;
      RECT  76.8 331.8 78.0 333.2 ;
      RECT  62.6 330.0 84.4 331.2 ;
      RECT  83.0 348.4 83.8 350.0 ;
      RECT  64.6 337.4 75.6 338.0 ;
      RECT  78.4 336.2 82.2 336.8 ;
      RECT  67.0 333.8 67.8 334.6 ;
      RECT  72.6 333.8 73.2 334.4 ;
      RECT  76.6 333.8 77.4 334.6 ;
      RECT  78.0 340.0 78.8 340.2 ;
      RECT  63.8 360.4 73.6 360.2 ;
      RECT  78.0 361.0 82.2 360.4 ;
      RECT  81.4 369.4 82.2 365.0 ;
      RECT  70.4 357.0 74.0 356.4 ;
      RECT  81.4 364.4 82.2 361.0 ;
      RECT  70.4 366.2 71.2 366.0 ;
      RECT  73.0 358.6 75.2 358.0 ;
      RECT  63.8 369.4 64.6 364.6 ;
      RECT  74.4 364.0 75.2 363.8 ;
      RECT  70.4 357.2 71.2 357.0 ;
      RECT  67.0 358.6 67.8 358.4 ;
      RECT  74.4 358.8 75.2 358.6 ;
      RECT  75.0 360.0 77.4 359.4 ;
      RECT  67.6 363.2 68.4 363.0 ;
      RECT  81.4 360.4 82.2 351.8 ;
      RECT  78.4 365.2 79.2 365.0 ;
      RECT  76.6 362.4 80.4 361.8 ;
      RECT  68.8 366.0 69.4 363.8 ;
      RECT  70.8 370.0 71.8 367.4 ;
      RECT  79.8 370.0 80.6 365.6 ;
      RECT  71.6 358.6 72.4 358.4 ;
      RECT  79.6 361.8 80.4 361.6 ;
      RECT  72.6 355.8 73.4 351.8 ;
      RECT  67.0 356.6 67.8 355.8 ;
      RECT  76.6 356.6 77.4 355.8 ;
      RECT  68.8 360.2 73.6 359.8 ;
      RECT  63.8 360.6 69.6 360.4 ;
      RECT  66.0 362.0 71.0 361.4 ;
      RECT  73.2 357.2 74.0 357.0 ;
      RECT  67.0 355.8 69.0 355.2 ;
      RECT  65.4 370.0 66.2 365.4 ;
      RECT  70.4 366.8 73.2 366.2 ;
      RECT  83.0 370.0 83.8 368.6 ;
      RECT  63.8 360.2 64.6 351.8 ;
      RECT  65.4 359.6 66.2 351.2 ;
      RECT  76.8 359.4 77.4 358.4 ;
      RECT  76.6 368.0 78.0 367.4 ;
      RECT  71.0 355.8 71.8 351.2 ;
      RECT  74.2 355.8 75.0 351.2 ;
      RECT  76.8 358.4 78.2 357.6 ;
      RECT  75.0 363.2 75.6 360.0 ;
      RECT  64.6 364.0 66.2 363.8 ;
      RECT  67.0 368.0 69.0 367.4 ;
      RECT  68.2 369.4 69.0 368.0 ;
      RECT  76.8 355.8 78.0 351.8 ;
      RECT  68.6 366.8 69.4 366.0 ;
      RECT  73.0 359.8 73.6 358.6 ;
      RECT  70.2 361.4 71.0 361.2 ;
      RECT  76.6 362.6 77.4 362.4 ;
      RECT  72.6 356.4 73.2 355.8 ;
      RECT  67.0 359.2 72.4 358.6 ;
      RECT  72.6 369.4 73.4 367.4 ;
      RECT  62.6 351.2 84.4 350.0 ;
      RECT  68.2 355.2 69.0 351.8 ;
      RECT  79.8 359.8 80.6 351.2 ;
      RECT  63.8 360.8 69.4 360.6 ;
      RECT  66.0 362.2 66.8 362.0 ;
      RECT  74.2 370.0 75.0 367.4 ;
      RECT  76.8 369.4 78.0 368.0 ;
      RECT  62.6 371.2 84.4 370.0 ;
      RECT  83.0 352.8 83.8 351.2 ;
      RECT  64.6 363.8 75.6 363.2 ;
      RECT  78.4 365.0 82.2 364.4 ;
      RECT  67.0 367.4 67.8 366.6 ;
      RECT  72.6 367.4 73.2 366.8 ;
      RECT  76.6 367.4 77.4 366.6 ;
      RECT  78.0 361.2 78.8 361.0 ;
      RECT  179.4 56.0 189.2 56.2 ;
      RECT  193.6 55.4 197.8 56.0 ;
      RECT  197.0 47.0 197.8 51.4 ;
      RECT  186.0 59.4 189.6 60.0 ;
      RECT  197.0 52.0 197.8 55.4 ;
      RECT  186.0 50.2 186.8 50.4 ;
      RECT  188.6 57.8 190.8 58.4 ;
      RECT  179.4 47.0 180.2 51.8 ;
      RECT  190.0 52.4 190.8 52.6 ;
      RECT  186.0 59.2 186.8 59.4 ;
      RECT  182.6 57.8 183.4 58.0 ;
      RECT  190.0 57.6 190.8 57.8 ;
      RECT  190.6 56.4 193.0 57.0 ;
      RECT  183.2 53.2 184.0 53.4 ;
      RECT  197.0 56.0 197.8 64.6 ;
      RECT  194.0 51.2 194.8 51.4 ;
      RECT  192.2 54.0 196.0 54.6 ;
      RECT  184.4 50.4 185.0 52.6 ;
      RECT  186.4 46.4 187.4 49.0 ;
      RECT  195.4 46.4 196.2 50.8 ;
      RECT  187.2 57.8 188.0 58.0 ;
      RECT  195.2 54.6 196.0 54.8 ;
      RECT  188.2 60.6 189.0 64.6 ;
      RECT  182.6 59.8 183.4 60.6 ;
      RECT  192.2 59.8 193.0 60.6 ;
      RECT  184.4 56.2 189.2 56.6 ;
      RECT  179.4 55.8 185.2 56.0 ;
      RECT  181.6 54.4 186.6 55.0 ;
      RECT  188.8 59.2 189.6 59.4 ;
      RECT  182.6 60.6 184.6 61.2 ;
      RECT  181.0 46.4 181.8 51.0 ;
      RECT  186.0 49.6 188.8 50.2 ;
      RECT  198.6 46.4 199.4 47.8 ;
      RECT  179.4 56.2 180.2 64.6 ;
      RECT  181.0 56.8 181.8 65.2 ;
      RECT  192.4 57.0 193.0 58.0 ;
      RECT  192.2 48.4 193.6 49.0 ;
      RECT  186.6 60.6 187.4 65.2 ;
      RECT  189.8 60.6 190.6 65.2 ;
      RECT  192.4 58.0 193.8 58.8 ;
      RECT  190.6 53.2 191.2 56.4 ;
      RECT  180.2 52.4 181.8 52.6 ;
      RECT  182.6 48.4 184.6 49.0 ;
      RECT  183.8 47.0 184.6 48.4 ;
      RECT  192.4 60.6 193.6 64.6 ;
      RECT  184.2 49.6 185.0 50.4 ;
      RECT  188.6 56.6 189.2 57.8 ;
      RECT  185.8 55.0 186.6 55.2 ;
      RECT  192.2 53.8 193.0 54.0 ;
      RECT  188.2 60.0 188.8 60.6 ;
      RECT  182.6 57.2 188.0 57.8 ;
      RECT  188.2 47.0 189.0 49.0 ;
      RECT  178.2 65.2 200.0 66.4 ;
      RECT  183.8 61.2 184.6 64.6 ;
      RECT  195.4 56.6 196.2 65.2 ;
      RECT  179.4 55.6 185.0 55.8 ;
      RECT  181.6 54.2 182.4 54.4 ;
      RECT  189.8 46.4 190.6 49.0 ;
      RECT  192.4 47.0 193.6 48.4 ;
      RECT  178.2 45.2 200.0 46.4 ;
      RECT  198.6 63.6 199.4 65.2 ;
      RECT  180.2 52.6 191.2 53.2 ;
      RECT  194.0 51.4 197.8 52.0 ;
      RECT  182.6 49.0 183.4 49.8 ;
      RECT  188.2 49.0 188.8 49.6 ;
      RECT  192.2 49.0 193.0 49.8 ;
      RECT  193.6 55.2 194.4 55.4 ;
      RECT  201.2 56.0 211.0 56.2 ;
      RECT  215.4 55.4 219.6 56.0 ;
      RECT  218.8 47.0 219.6 51.4 ;
      RECT  207.8 59.4 211.4 60.0 ;
      RECT  218.8 52.0 219.6 55.4 ;
      RECT  207.8 50.2 208.6 50.4 ;
      RECT  210.4 57.8 212.6 58.4 ;
      RECT  201.2 47.0 202.0 51.8 ;
      RECT  211.8 52.4 212.6 52.6 ;
      RECT  207.8 59.2 208.6 59.4 ;
      RECT  204.4 57.8 205.2 58.0 ;
      RECT  211.8 57.6 212.6 57.8 ;
      RECT  212.4 56.4 214.8 57.0 ;
      RECT  205.0 53.2 205.8 53.4 ;
      RECT  218.8 56.0 219.6 64.6 ;
      RECT  215.8 51.2 216.6 51.4 ;
      RECT  214.0 54.0 217.8 54.6 ;
      RECT  206.2 50.4 206.8 52.6 ;
      RECT  208.2 46.4 209.2 49.0 ;
      RECT  217.2 46.4 218.0 50.8 ;
      RECT  209.0 57.8 209.8 58.0 ;
      RECT  217.0 54.6 217.8 54.8 ;
      RECT  210.0 60.6 210.8 64.6 ;
      RECT  204.4 59.8 205.2 60.6 ;
      RECT  214.0 59.8 214.8 60.6 ;
      RECT  206.2 56.2 211.0 56.6 ;
      RECT  201.2 55.8 207.0 56.0 ;
      RECT  203.4 54.4 208.4 55.0 ;
      RECT  210.6 59.2 211.4 59.4 ;
      RECT  204.4 60.6 206.4 61.2 ;
      RECT  202.8 46.4 203.6 51.0 ;
      RECT  207.8 49.6 210.6 50.2 ;
      RECT  220.4 46.4 221.2 47.8 ;
      RECT  201.2 56.2 202.0 64.6 ;
      RECT  202.8 56.8 203.6 65.2 ;
      RECT  214.2 57.0 214.8 58.0 ;
      RECT  214.0 48.4 215.4 49.0 ;
      RECT  208.4 60.6 209.2 65.2 ;
      RECT  211.6 60.6 212.4 65.2 ;
      RECT  214.2 58.0 215.6 58.8 ;
      RECT  212.4 53.2 213.0 56.4 ;
      RECT  202.0 52.4 203.6 52.6 ;
      RECT  204.4 48.4 206.4 49.0 ;
      RECT  205.6 47.0 206.4 48.4 ;
      RECT  214.2 60.6 215.4 64.6 ;
      RECT  206.0 49.6 206.8 50.4 ;
      RECT  210.4 56.6 211.0 57.8 ;
      RECT  207.6 55.0 208.4 55.2 ;
      RECT  214.0 53.8 214.8 54.0 ;
      RECT  210.0 60.0 210.6 60.6 ;
      RECT  204.4 57.2 209.8 57.8 ;
      RECT  210.0 47.0 210.8 49.0 ;
      RECT  200.0 65.2 221.8 66.4 ;
      RECT  205.6 61.2 206.4 64.6 ;
      RECT  217.2 56.6 218.0 65.2 ;
      RECT  201.2 55.6 206.8 55.8 ;
      RECT  203.4 54.2 204.2 54.4 ;
      RECT  211.6 46.4 212.4 49.0 ;
      RECT  214.2 47.0 215.4 48.4 ;
      RECT  200.0 45.2 221.8 46.4 ;
      RECT  220.4 63.6 221.2 65.2 ;
      RECT  202.0 52.6 213.0 53.2 ;
      RECT  215.8 51.4 219.6 52.0 ;
      RECT  204.4 49.0 205.2 49.8 ;
      RECT  210.0 49.0 210.6 49.6 ;
      RECT  214.0 49.0 214.8 49.8 ;
      RECT  215.4 55.2 216.2 55.4 ;
   LAYER  m2 ;
      RECT  191.4 192.0 192.2 202.8 ;
      RECT  194.8 202.0 195.6 202.8 ;
      RECT  196.6 193.6 197.4 202.8 ;
      RECT  193.0 192.0 193.8 202.8 ;
      RECT  198.2 192.0 199.0 202.8 ;
      RECT  195.8 192.8 197.4 193.6 ;
      RECT  196.6 192.0 197.4 192.8 ;
      RECT  191.4 212.8 192.2 202.0 ;
      RECT  194.8 202.8 195.6 202.0 ;
      RECT  196.6 211.2 197.4 202.0 ;
      RECT  193.0 212.8 193.8 202.0 ;
      RECT  198.2 212.8 199.0 202.0 ;
      RECT  195.8 212.0 197.4 211.2 ;
      RECT  196.6 212.8 197.4 212.0 ;
      RECT  191.4 212.8 192.2 223.6 ;
      RECT  194.8 222.8 195.6 223.6 ;
      RECT  196.6 214.4 197.4 223.6 ;
      RECT  193.0 212.8 193.8 223.6 ;
      RECT  198.2 212.8 199.0 223.6 ;
      RECT  195.8 213.6 197.4 214.4 ;
      RECT  196.6 212.8 197.4 213.6 ;
      RECT  191.4 233.6 192.2 222.8 ;
      RECT  194.8 223.6 195.6 222.8 ;
      RECT  196.6 232.0 197.4 222.8 ;
      RECT  193.0 233.6 193.8 222.8 ;
      RECT  198.2 233.6 199.0 222.8 ;
      RECT  195.8 232.8 197.4 232.0 ;
      RECT  196.6 233.6 197.4 232.8 ;
      RECT  191.4 233.6 192.2 244.4 ;
      RECT  194.8 243.6 195.6 244.4 ;
      RECT  196.6 235.2 197.4 244.4 ;
      RECT  193.0 233.6 193.8 244.4 ;
      RECT  198.2 233.6 199.0 244.4 ;
      RECT  195.8 234.4 197.4 235.2 ;
      RECT  196.6 233.6 197.4 234.4 ;
      RECT  191.4 254.4 192.2 243.6 ;
      RECT  194.8 244.4 195.6 243.6 ;
      RECT  196.6 252.8 197.4 243.6 ;
      RECT  193.0 254.4 193.8 243.6 ;
      RECT  198.2 254.4 199.0 243.6 ;
      RECT  195.8 253.6 197.4 252.8 ;
      RECT  196.6 254.4 197.4 253.6 ;
      RECT  191.4 254.4 192.2 265.2 ;
      RECT  194.8 264.4 195.6 265.2 ;
      RECT  196.6 256.0 197.4 265.2 ;
      RECT  193.0 254.4 193.8 265.2 ;
      RECT  198.2 254.4 199.0 265.2 ;
      RECT  195.8 255.2 197.4 256.0 ;
      RECT  196.6 254.4 197.4 255.2 ;
      RECT  191.4 275.2 192.2 264.4 ;
      RECT  194.8 265.2 195.6 264.4 ;
      RECT  196.6 273.6 197.4 264.4 ;
      RECT  193.0 275.2 193.8 264.4 ;
      RECT  198.2 275.2 199.0 264.4 ;
      RECT  195.8 274.4 197.4 273.6 ;
      RECT  196.6 275.2 197.4 274.4 ;
      RECT  191.4 275.2 192.2 286.0 ;
      RECT  194.8 285.2 195.6 286.0 ;
      RECT  196.6 276.8 197.4 286.0 ;
      RECT  193.0 275.2 193.8 286.0 ;
      RECT  198.2 275.2 199.0 286.0 ;
      RECT  195.8 276.0 197.4 276.8 ;
      RECT  196.6 275.2 197.4 276.0 ;
      RECT  191.4 296.0 192.2 285.2 ;
      RECT  194.8 286.0 195.6 285.2 ;
      RECT  196.6 294.4 197.4 285.2 ;
      RECT  193.0 296.0 193.8 285.2 ;
      RECT  198.2 296.0 199.0 285.2 ;
      RECT  195.8 295.2 197.4 294.4 ;
      RECT  196.6 296.0 197.4 295.2 ;
      RECT  191.4 296.0 192.2 306.8 ;
      RECT  194.8 306.0 195.6 306.8 ;
      RECT  196.6 297.6 197.4 306.8 ;
      RECT  193.0 296.0 193.8 306.8 ;
      RECT  198.2 296.0 199.0 306.8 ;
      RECT  195.8 296.8 197.4 297.6 ;
      RECT  196.6 296.0 197.4 296.8 ;
      RECT  191.4 316.8 192.2 306.0 ;
      RECT  194.8 306.8 195.6 306.0 ;
      RECT  196.6 315.2 197.4 306.0 ;
      RECT  193.0 316.8 193.8 306.0 ;
      RECT  198.2 316.8 199.0 306.0 ;
      RECT  195.8 316.0 197.4 315.2 ;
      RECT  196.6 316.8 197.4 316.0 ;
      RECT  191.4 316.8 192.2 327.6 ;
      RECT  194.8 326.8 195.6 327.6 ;
      RECT  196.6 318.4 197.4 327.6 ;
      RECT  193.0 316.8 193.8 327.6 ;
      RECT  198.2 316.8 199.0 327.6 ;
      RECT  195.8 317.6 197.4 318.4 ;
      RECT  196.6 316.8 197.4 317.6 ;
      RECT  191.4 337.6 192.2 326.8 ;
      RECT  194.8 327.6 195.6 326.8 ;
      RECT  196.6 336.0 197.4 326.8 ;
      RECT  193.0 337.6 193.8 326.8 ;
      RECT  198.2 337.6 199.0 326.8 ;
      RECT  195.8 336.8 197.4 336.0 ;
      RECT  196.6 337.6 197.4 336.8 ;
      RECT  191.4 337.6 192.2 348.4 ;
      RECT  194.8 347.6 195.6 348.4 ;
      RECT  196.6 339.2 197.4 348.4 ;
      RECT  193.0 337.6 193.8 348.4 ;
      RECT  198.2 337.6 199.0 348.4 ;
      RECT  195.8 338.4 197.4 339.2 ;
      RECT  196.6 337.6 197.4 338.4 ;
      RECT  191.4 358.4 192.2 347.6 ;
      RECT  194.8 348.4 195.6 347.6 ;
      RECT  196.6 356.8 197.4 347.6 ;
      RECT  193.0 358.4 193.8 347.6 ;
      RECT  198.2 358.4 199.0 347.6 ;
      RECT  195.8 357.6 197.4 356.8 ;
      RECT  196.6 358.4 197.4 357.6 ;
      RECT  198.2 192.0 199.0 202.8 ;
      RECT  201.6 202.0 202.4 202.8 ;
      RECT  203.4 193.6 204.2 202.8 ;
      RECT  199.8 192.0 200.6 202.8 ;
      RECT  205.0 192.0 205.8 202.8 ;
      RECT  202.6 192.8 204.2 193.6 ;
      RECT  203.4 192.0 204.2 192.8 ;
      RECT  198.2 212.8 199.0 202.0 ;
      RECT  201.6 202.8 202.4 202.0 ;
      RECT  203.4 211.2 204.2 202.0 ;
      RECT  199.8 212.8 200.6 202.0 ;
      RECT  205.0 212.8 205.8 202.0 ;
      RECT  202.6 212.0 204.2 211.2 ;
      RECT  203.4 212.8 204.2 212.0 ;
      RECT  198.2 212.8 199.0 223.6 ;
      RECT  201.6 222.8 202.4 223.6 ;
      RECT  203.4 214.4 204.2 223.6 ;
      RECT  199.8 212.8 200.6 223.6 ;
      RECT  205.0 212.8 205.8 223.6 ;
      RECT  202.6 213.6 204.2 214.4 ;
      RECT  203.4 212.8 204.2 213.6 ;
      RECT  198.2 233.6 199.0 222.8 ;
      RECT  201.6 223.6 202.4 222.8 ;
      RECT  203.4 232.0 204.2 222.8 ;
      RECT  199.8 233.6 200.6 222.8 ;
      RECT  205.0 233.6 205.8 222.8 ;
      RECT  202.6 232.8 204.2 232.0 ;
      RECT  203.4 233.6 204.2 232.8 ;
      RECT  198.2 233.6 199.0 244.4 ;
      RECT  201.6 243.6 202.4 244.4 ;
      RECT  203.4 235.2 204.2 244.4 ;
      RECT  199.8 233.6 200.6 244.4 ;
      RECT  205.0 233.6 205.8 244.4 ;
      RECT  202.6 234.4 204.2 235.2 ;
      RECT  203.4 233.6 204.2 234.4 ;
      RECT  198.2 254.4 199.0 243.6 ;
      RECT  201.6 244.4 202.4 243.6 ;
      RECT  203.4 252.8 204.2 243.6 ;
      RECT  199.8 254.4 200.6 243.6 ;
      RECT  205.0 254.4 205.8 243.6 ;
      RECT  202.6 253.6 204.2 252.8 ;
      RECT  203.4 254.4 204.2 253.6 ;
      RECT  198.2 254.4 199.0 265.2 ;
      RECT  201.6 264.4 202.4 265.2 ;
      RECT  203.4 256.0 204.2 265.2 ;
      RECT  199.8 254.4 200.6 265.2 ;
      RECT  205.0 254.4 205.8 265.2 ;
      RECT  202.6 255.2 204.2 256.0 ;
      RECT  203.4 254.4 204.2 255.2 ;
      RECT  198.2 275.2 199.0 264.4 ;
      RECT  201.6 265.2 202.4 264.4 ;
      RECT  203.4 273.6 204.2 264.4 ;
      RECT  199.8 275.2 200.6 264.4 ;
      RECT  205.0 275.2 205.8 264.4 ;
      RECT  202.6 274.4 204.2 273.6 ;
      RECT  203.4 275.2 204.2 274.4 ;
      RECT  198.2 275.2 199.0 286.0 ;
      RECT  201.6 285.2 202.4 286.0 ;
      RECT  203.4 276.8 204.2 286.0 ;
      RECT  199.8 275.2 200.6 286.0 ;
      RECT  205.0 275.2 205.8 286.0 ;
      RECT  202.6 276.0 204.2 276.8 ;
      RECT  203.4 275.2 204.2 276.0 ;
      RECT  198.2 296.0 199.0 285.2 ;
      RECT  201.6 286.0 202.4 285.2 ;
      RECT  203.4 294.4 204.2 285.2 ;
      RECT  199.8 296.0 200.6 285.2 ;
      RECT  205.0 296.0 205.8 285.2 ;
      RECT  202.6 295.2 204.2 294.4 ;
      RECT  203.4 296.0 204.2 295.2 ;
      RECT  198.2 296.0 199.0 306.8 ;
      RECT  201.6 306.0 202.4 306.8 ;
      RECT  203.4 297.6 204.2 306.8 ;
      RECT  199.8 296.0 200.6 306.8 ;
      RECT  205.0 296.0 205.8 306.8 ;
      RECT  202.6 296.8 204.2 297.6 ;
      RECT  203.4 296.0 204.2 296.8 ;
      RECT  198.2 316.8 199.0 306.0 ;
      RECT  201.6 306.8 202.4 306.0 ;
      RECT  203.4 315.2 204.2 306.0 ;
      RECT  199.8 316.8 200.6 306.0 ;
      RECT  205.0 316.8 205.8 306.0 ;
      RECT  202.6 316.0 204.2 315.2 ;
      RECT  203.4 316.8 204.2 316.0 ;
      RECT  198.2 316.8 199.0 327.6 ;
      RECT  201.6 326.8 202.4 327.6 ;
      RECT  203.4 318.4 204.2 327.6 ;
      RECT  199.8 316.8 200.6 327.6 ;
      RECT  205.0 316.8 205.8 327.6 ;
      RECT  202.6 317.6 204.2 318.4 ;
      RECT  203.4 316.8 204.2 317.6 ;
      RECT  198.2 337.6 199.0 326.8 ;
      RECT  201.6 327.6 202.4 326.8 ;
      RECT  203.4 336.0 204.2 326.8 ;
      RECT  199.8 337.6 200.6 326.8 ;
      RECT  205.0 337.6 205.8 326.8 ;
      RECT  202.6 336.8 204.2 336.0 ;
      RECT  203.4 337.6 204.2 336.8 ;
      RECT  198.2 337.6 199.0 348.4 ;
      RECT  201.6 347.6 202.4 348.4 ;
      RECT  203.4 339.2 204.2 348.4 ;
      RECT  199.8 337.6 200.6 348.4 ;
      RECT  205.0 337.6 205.8 348.4 ;
      RECT  202.6 338.4 204.2 339.2 ;
      RECT  203.4 337.6 204.2 338.4 ;
      RECT  198.2 358.4 199.0 347.6 ;
      RECT  201.6 348.4 202.4 347.6 ;
      RECT  203.4 356.8 204.2 347.6 ;
      RECT  199.8 358.4 200.6 347.6 ;
      RECT  205.0 358.4 205.8 347.6 ;
      RECT  202.6 357.6 204.2 356.8 ;
      RECT  203.4 358.4 204.2 357.6 ;
      RECT  193.0 192.0 193.8 358.4 ;
      RECT  196.6 192.0 197.4 358.4 ;
      RECT  199.8 192.0 200.6 358.4 ;
      RECT  203.4 192.0 204.2 358.4 ;
      RECT  191.4 171.2 192.2 182.0 ;
      RECT  184.6 171.2 185.4 182.0 ;
      RECT  188.0 181.2 188.8 182.0 ;
      RECT  189.8 171.2 190.6 182.0 ;
      RECT  186.2 171.2 187.0 182.0 ;
      RECT  184.6 192.0 185.4 181.2 ;
      RECT  188.0 182.0 188.8 181.2 ;
      RECT  189.8 190.4 190.6 181.2 ;
      RECT  186.2 192.0 187.0 181.2 ;
      RECT  191.4 192.0 192.2 181.2 ;
      RECT  189.0 191.2 190.6 190.4 ;
      RECT  189.8 192.0 190.6 191.2 ;
      RECT  184.6 192.0 185.4 202.8 ;
      RECT  188.0 202.0 188.8 202.8 ;
      RECT  189.8 193.6 190.6 202.8 ;
      RECT  186.2 192.0 187.0 202.8 ;
      RECT  191.4 192.0 192.2 202.8 ;
      RECT  189.0 192.8 190.6 193.6 ;
      RECT  189.8 192.0 190.6 192.8 ;
      RECT  184.6 212.8 185.4 202.0 ;
      RECT  188.0 202.8 188.8 202.0 ;
      RECT  189.8 211.2 190.6 202.0 ;
      RECT  186.2 212.8 187.0 202.0 ;
      RECT  191.4 212.8 192.2 202.0 ;
      RECT  189.0 212.0 190.6 211.2 ;
      RECT  189.8 212.8 190.6 212.0 ;
      RECT  184.6 212.8 185.4 223.6 ;
      RECT  188.0 222.8 188.8 223.6 ;
      RECT  189.8 214.4 190.6 223.6 ;
      RECT  186.2 212.8 187.0 223.6 ;
      RECT  191.4 212.8 192.2 223.6 ;
      RECT  189.0 213.6 190.6 214.4 ;
      RECT  189.8 212.8 190.6 213.6 ;
      RECT  184.6 233.6 185.4 222.8 ;
      RECT  188.0 223.6 188.8 222.8 ;
      RECT  189.8 232.0 190.6 222.8 ;
      RECT  186.2 233.6 187.0 222.8 ;
      RECT  191.4 233.6 192.2 222.8 ;
      RECT  189.0 232.8 190.6 232.0 ;
      RECT  189.8 233.6 190.6 232.8 ;
      RECT  184.6 233.6 185.4 244.4 ;
      RECT  188.0 243.6 188.8 244.4 ;
      RECT  189.8 235.2 190.6 244.4 ;
      RECT  186.2 233.6 187.0 244.4 ;
      RECT  191.4 233.6 192.2 244.4 ;
      RECT  189.0 234.4 190.6 235.2 ;
      RECT  189.8 233.6 190.6 234.4 ;
      RECT  184.6 254.4 185.4 243.6 ;
      RECT  188.0 244.4 188.8 243.6 ;
      RECT  189.8 252.8 190.6 243.6 ;
      RECT  186.2 254.4 187.0 243.6 ;
      RECT  191.4 254.4 192.2 243.6 ;
      RECT  189.0 253.6 190.6 252.8 ;
      RECT  189.8 254.4 190.6 253.6 ;
      RECT  184.6 254.4 185.4 265.2 ;
      RECT  188.0 264.4 188.8 265.2 ;
      RECT  189.8 256.0 190.6 265.2 ;
      RECT  186.2 254.4 187.0 265.2 ;
      RECT  191.4 254.4 192.2 265.2 ;
      RECT  189.0 255.2 190.6 256.0 ;
      RECT  189.8 254.4 190.6 255.2 ;
      RECT  184.6 275.2 185.4 264.4 ;
      RECT  188.0 265.2 188.8 264.4 ;
      RECT  189.8 273.6 190.6 264.4 ;
      RECT  186.2 275.2 187.0 264.4 ;
      RECT  191.4 275.2 192.2 264.4 ;
      RECT  189.0 274.4 190.6 273.6 ;
      RECT  189.8 275.2 190.6 274.4 ;
      RECT  184.6 275.2 185.4 286.0 ;
      RECT  188.0 285.2 188.8 286.0 ;
      RECT  189.8 276.8 190.6 286.0 ;
      RECT  186.2 275.2 187.0 286.0 ;
      RECT  191.4 275.2 192.2 286.0 ;
      RECT  189.0 276.0 190.6 276.8 ;
      RECT  189.8 275.2 190.6 276.0 ;
      RECT  184.6 296.0 185.4 285.2 ;
      RECT  188.0 286.0 188.8 285.2 ;
      RECT  189.8 294.4 190.6 285.2 ;
      RECT  186.2 296.0 187.0 285.2 ;
      RECT  191.4 296.0 192.2 285.2 ;
      RECT  189.0 295.2 190.6 294.4 ;
      RECT  189.8 296.0 190.6 295.2 ;
      RECT  184.6 296.0 185.4 306.8 ;
      RECT  188.0 306.0 188.8 306.8 ;
      RECT  189.8 297.6 190.6 306.8 ;
      RECT  186.2 296.0 187.0 306.8 ;
      RECT  191.4 296.0 192.2 306.8 ;
      RECT  189.0 296.8 190.6 297.6 ;
      RECT  189.8 296.0 190.6 296.8 ;
      RECT  184.6 316.8 185.4 306.0 ;
      RECT  188.0 306.8 188.8 306.0 ;
      RECT  189.8 315.2 190.6 306.0 ;
      RECT  186.2 316.8 187.0 306.0 ;
      RECT  191.4 316.8 192.2 306.0 ;
      RECT  189.0 316.0 190.6 315.2 ;
      RECT  189.8 316.8 190.6 316.0 ;
      RECT  184.6 316.8 185.4 327.6 ;
      RECT  188.0 326.8 188.8 327.6 ;
      RECT  189.8 318.4 190.6 327.6 ;
      RECT  186.2 316.8 187.0 327.6 ;
      RECT  191.4 316.8 192.2 327.6 ;
      RECT  189.0 317.6 190.6 318.4 ;
      RECT  189.8 316.8 190.6 317.6 ;
      RECT  184.6 337.6 185.4 326.8 ;
      RECT  188.0 327.6 188.8 326.8 ;
      RECT  189.8 336.0 190.6 326.8 ;
      RECT  186.2 337.6 187.0 326.8 ;
      RECT  191.4 337.6 192.2 326.8 ;
      RECT  189.0 336.8 190.6 336.0 ;
      RECT  189.8 337.6 190.6 336.8 ;
      RECT  184.6 337.6 185.4 348.4 ;
      RECT  188.0 347.6 188.8 348.4 ;
      RECT  189.8 339.2 190.6 348.4 ;
      RECT  186.2 337.6 187.0 348.4 ;
      RECT  191.4 337.6 192.2 348.4 ;
      RECT  189.0 338.4 190.6 339.2 ;
      RECT  189.8 337.6 190.6 338.4 ;
      RECT  184.6 358.4 185.4 347.6 ;
      RECT  188.0 348.4 188.8 347.6 ;
      RECT  189.8 356.8 190.6 347.6 ;
      RECT  186.2 358.4 187.0 347.6 ;
      RECT  191.4 358.4 192.2 347.6 ;
      RECT  189.0 357.6 190.6 356.8 ;
      RECT  189.8 358.4 190.6 357.6 ;
      RECT  191.4 358.4 192.2 369.2 ;
      RECT  184.6 358.4 185.4 369.2 ;
      RECT  188.0 368.4 188.8 369.2 ;
      RECT  189.8 358.4 190.6 369.2 ;
      RECT  186.2 358.4 187.0 369.2 ;
      RECT  188.0 326.8 188.8 327.6 ;
      RECT  188.0 264.4 188.8 265.2 ;
      RECT  188.0 202.0 188.8 202.8 ;
      RECT  188.0 285.2 188.8 286.0 ;
      RECT  188.0 285.2 188.8 286.0 ;
      RECT  188.0 181.2 188.8 182.0 ;
      RECT  188.0 306.0 188.8 306.8 ;
      RECT  188.0 306.0 188.8 306.8 ;
      RECT  188.0 222.8 188.8 223.6 ;
      RECT  188.0 222.8 188.8 223.6 ;
      RECT  188.0 243.6 188.8 244.4 ;
      RECT  188.0 368.4 188.8 369.2 ;
      RECT  188.0 347.6 188.8 348.4 ;
      RECT  184.6 212.8 185.4 223.6 ;
      RECT  191.4 181.2 192.2 192.0 ;
      RECT  184.6 285.2 185.4 296.0 ;
      RECT  191.4 285.2 192.2 296.0 ;
      RECT  184.6 306.0 185.4 316.8 ;
      RECT  184.6 202.0 185.4 212.8 ;
      RECT  184.6 275.2 185.4 286.0 ;
      RECT  184.6 316.8 185.4 327.6 ;
      RECT  184.6 337.6 185.4 348.4 ;
      RECT  184.6 358.4 185.4 369.2 ;
      RECT  191.4 275.2 192.2 286.0 ;
      RECT  191.4 233.6 192.2 244.4 ;
      RECT  191.4 358.4 192.2 369.2 ;
      RECT  191.4 171.2 192.2 182.0 ;
      RECT  184.6 243.6 185.4 254.4 ;
      RECT  191.4 296.0 192.2 306.8 ;
      RECT  191.4 264.4 192.2 275.2 ;
      RECT  184.6 181.2 185.4 192.0 ;
      RECT  191.4 337.6 192.2 348.4 ;
      RECT  191.4 306.0 192.2 316.8 ;
      RECT  191.4 212.8 192.2 223.6 ;
      RECT  184.6 347.6 185.4 358.4 ;
      RECT  184.6 192.0 185.4 202.8 ;
      RECT  184.6 264.4 185.4 275.2 ;
      RECT  184.6 326.8 185.4 337.6 ;
      RECT  191.4 192.0 192.2 202.8 ;
      RECT  184.6 171.2 185.4 182.0 ;
      RECT  184.6 222.8 185.4 233.6 ;
      RECT  191.4 254.4 192.2 265.2 ;
      RECT  191.4 202.0 192.2 212.8 ;
      RECT  184.6 296.0 185.4 306.8 ;
      RECT  191.4 326.8 192.2 337.6 ;
      RECT  191.4 347.6 192.2 358.4 ;
      RECT  184.6 254.4 185.4 265.2 ;
      RECT  184.6 233.6 185.4 244.4 ;
      RECT  191.4 222.8 192.2 233.6 ;
      RECT  191.4 316.8 192.2 327.6 ;
      RECT  191.4 243.6 192.2 254.4 ;
      RECT  198.2 192.0 199.0 181.2 ;
      RECT  191.4 192.0 192.2 181.2 ;
      RECT  194.8 182.0 195.6 181.2 ;
      RECT  196.6 192.0 197.4 181.2 ;
      RECT  193.0 192.0 193.8 181.2 ;
      RECT  205.0 192.0 205.8 181.2 ;
      RECT  198.2 192.0 199.0 181.2 ;
      RECT  201.6 182.0 202.4 181.2 ;
      RECT  203.4 192.0 204.2 181.2 ;
      RECT  199.8 192.0 200.6 181.2 ;
      RECT  193.0 192.0 193.8 181.6 ;
      RECT  196.6 192.0 197.4 181.6 ;
      RECT  199.8 192.0 200.6 181.6 ;
      RECT  203.4 192.0 204.2 181.6 ;
      RECT  198.2 171.2 199.0 182.0 ;
      RECT  191.4 171.2 192.2 182.0 ;
      RECT  194.8 181.2 195.6 182.0 ;
      RECT  196.6 171.2 197.4 182.0 ;
      RECT  193.0 171.2 193.8 182.0 ;
      RECT  205.0 171.2 205.8 182.0 ;
      RECT  198.2 171.2 199.0 182.0 ;
      RECT  201.6 181.2 202.4 182.0 ;
      RECT  203.4 171.2 204.2 182.0 ;
      RECT  199.8 171.2 200.6 182.0 ;
      RECT  193.0 171.2 193.8 181.6 ;
      RECT  196.6 171.2 197.4 181.6 ;
      RECT  199.8 171.2 200.6 181.6 ;
      RECT  203.4 171.2 204.2 181.6 ;
      RECT  198.2 358.4 199.0 369.2 ;
      RECT  191.4 358.4 192.2 369.2 ;
      RECT  194.8 368.4 195.6 369.2 ;
      RECT  196.6 358.4 197.4 369.2 ;
      RECT  193.0 358.4 193.8 369.2 ;
      RECT  205.0 358.4 205.8 369.2 ;
      RECT  198.2 358.4 199.0 369.2 ;
      RECT  201.6 368.4 202.4 369.2 ;
      RECT  203.4 358.4 204.2 369.2 ;
      RECT  199.8 358.4 200.6 369.2 ;
      RECT  193.0 358.4 193.8 368.8 ;
      RECT  196.6 358.4 197.4 368.8 ;
      RECT  199.8 358.4 200.6 368.8 ;
      RECT  203.4 358.4 204.2 368.8 ;
      RECT  184.6 171.2 185.4 182.0 ;
      RECT  177.8 171.2 178.6 182.0 ;
      RECT  181.2 181.2 182.0 182.0 ;
      RECT  183.0 171.2 183.8 182.0 ;
      RECT  179.4 171.2 180.2 182.0 ;
      RECT  184.6 192.0 185.4 181.2 ;
      RECT  177.8 192.0 178.6 181.2 ;
      RECT  181.2 182.0 182.0 181.2 ;
      RECT  183.0 192.0 183.8 181.2 ;
      RECT  179.4 192.0 180.2 181.2 ;
      RECT  184.6 192.0 185.4 202.8 ;
      RECT  177.8 192.0 178.6 202.8 ;
      RECT  181.2 202.0 182.0 202.8 ;
      RECT  183.0 192.0 183.8 202.8 ;
      RECT  179.4 192.0 180.2 202.8 ;
      RECT  184.6 212.8 185.4 202.0 ;
      RECT  177.8 212.8 178.6 202.0 ;
      RECT  181.2 202.8 182.0 202.0 ;
      RECT  183.0 212.8 183.8 202.0 ;
      RECT  179.4 212.8 180.2 202.0 ;
      RECT  184.6 212.8 185.4 223.6 ;
      RECT  177.8 212.8 178.6 223.6 ;
      RECT  181.2 222.8 182.0 223.6 ;
      RECT  183.0 212.8 183.8 223.6 ;
      RECT  179.4 212.8 180.2 223.6 ;
      RECT  184.6 233.6 185.4 222.8 ;
      RECT  177.8 233.6 178.6 222.8 ;
      RECT  181.2 223.6 182.0 222.8 ;
      RECT  183.0 233.6 183.8 222.8 ;
      RECT  179.4 233.6 180.2 222.8 ;
      RECT  184.6 233.6 185.4 244.4 ;
      RECT  177.8 233.6 178.6 244.4 ;
      RECT  181.2 243.6 182.0 244.4 ;
      RECT  183.0 233.6 183.8 244.4 ;
      RECT  179.4 233.6 180.2 244.4 ;
      RECT  184.6 254.4 185.4 243.6 ;
      RECT  177.8 254.4 178.6 243.6 ;
      RECT  181.2 244.4 182.0 243.6 ;
      RECT  183.0 254.4 183.8 243.6 ;
      RECT  179.4 254.4 180.2 243.6 ;
      RECT  184.6 254.4 185.4 265.2 ;
      RECT  177.8 254.4 178.6 265.2 ;
      RECT  181.2 264.4 182.0 265.2 ;
      RECT  183.0 254.4 183.8 265.2 ;
      RECT  179.4 254.4 180.2 265.2 ;
      RECT  184.6 275.2 185.4 264.4 ;
      RECT  177.8 275.2 178.6 264.4 ;
      RECT  181.2 265.2 182.0 264.4 ;
      RECT  183.0 275.2 183.8 264.4 ;
      RECT  179.4 275.2 180.2 264.4 ;
      RECT  184.6 275.2 185.4 286.0 ;
      RECT  177.8 275.2 178.6 286.0 ;
      RECT  181.2 285.2 182.0 286.0 ;
      RECT  183.0 275.2 183.8 286.0 ;
      RECT  179.4 275.2 180.2 286.0 ;
      RECT  184.6 296.0 185.4 285.2 ;
      RECT  177.8 296.0 178.6 285.2 ;
      RECT  181.2 286.0 182.0 285.2 ;
      RECT  183.0 296.0 183.8 285.2 ;
      RECT  179.4 296.0 180.2 285.2 ;
      RECT  184.6 296.0 185.4 306.8 ;
      RECT  177.8 296.0 178.6 306.8 ;
      RECT  181.2 306.0 182.0 306.8 ;
      RECT  183.0 296.0 183.8 306.8 ;
      RECT  179.4 296.0 180.2 306.8 ;
      RECT  184.6 316.8 185.4 306.0 ;
      RECT  177.8 316.8 178.6 306.0 ;
      RECT  181.2 306.8 182.0 306.0 ;
      RECT  183.0 316.8 183.8 306.0 ;
      RECT  179.4 316.8 180.2 306.0 ;
      RECT  184.6 316.8 185.4 327.6 ;
      RECT  177.8 316.8 178.6 327.6 ;
      RECT  181.2 326.8 182.0 327.6 ;
      RECT  183.0 316.8 183.8 327.6 ;
      RECT  179.4 316.8 180.2 327.6 ;
      RECT  184.6 337.6 185.4 326.8 ;
      RECT  177.8 337.6 178.6 326.8 ;
      RECT  181.2 327.6 182.0 326.8 ;
      RECT  183.0 337.6 183.8 326.8 ;
      RECT  179.4 337.6 180.2 326.8 ;
      RECT  184.6 337.6 185.4 348.4 ;
      RECT  177.8 337.6 178.6 348.4 ;
      RECT  181.2 347.6 182.0 348.4 ;
      RECT  183.0 337.6 183.8 348.4 ;
      RECT  179.4 337.6 180.2 348.4 ;
      RECT  184.6 358.4 185.4 347.6 ;
      RECT  177.8 358.4 178.6 347.6 ;
      RECT  181.2 348.4 182.0 347.6 ;
      RECT  183.0 358.4 183.8 347.6 ;
      RECT  179.4 358.4 180.2 347.6 ;
      RECT  184.6 358.4 185.4 369.2 ;
      RECT  177.8 358.4 178.6 369.2 ;
      RECT  181.2 368.4 182.0 369.2 ;
      RECT  183.0 358.4 183.8 369.2 ;
      RECT  179.4 358.4 180.2 369.2 ;
      RECT  179.4 171.2 180.2 368.8 ;
      RECT  183.0 171.2 183.8 368.8 ;
      RECT  211.8 171.2 212.6 182.0 ;
      RECT  205.0 171.2 205.8 182.0 ;
      RECT  208.4 181.2 209.2 182.0 ;
      RECT  210.2 171.2 211.0 182.0 ;
      RECT  206.6 171.2 207.4 182.0 ;
      RECT  211.8 192.0 212.6 181.2 ;
      RECT  205.0 192.0 205.8 181.2 ;
      RECT  208.4 182.0 209.2 181.2 ;
      RECT  210.2 192.0 211.0 181.2 ;
      RECT  206.6 192.0 207.4 181.2 ;
      RECT  211.8 192.0 212.6 202.8 ;
      RECT  205.0 192.0 205.8 202.8 ;
      RECT  208.4 202.0 209.2 202.8 ;
      RECT  210.2 192.0 211.0 202.8 ;
      RECT  206.6 192.0 207.4 202.8 ;
      RECT  211.8 212.8 212.6 202.0 ;
      RECT  205.0 212.8 205.8 202.0 ;
      RECT  208.4 202.8 209.2 202.0 ;
      RECT  210.2 212.8 211.0 202.0 ;
      RECT  206.6 212.8 207.4 202.0 ;
      RECT  211.8 212.8 212.6 223.6 ;
      RECT  205.0 212.8 205.8 223.6 ;
      RECT  208.4 222.8 209.2 223.6 ;
      RECT  210.2 212.8 211.0 223.6 ;
      RECT  206.6 212.8 207.4 223.6 ;
      RECT  211.8 233.6 212.6 222.8 ;
      RECT  205.0 233.6 205.8 222.8 ;
      RECT  208.4 223.6 209.2 222.8 ;
      RECT  210.2 233.6 211.0 222.8 ;
      RECT  206.6 233.6 207.4 222.8 ;
      RECT  211.8 233.6 212.6 244.4 ;
      RECT  205.0 233.6 205.8 244.4 ;
      RECT  208.4 243.6 209.2 244.4 ;
      RECT  210.2 233.6 211.0 244.4 ;
      RECT  206.6 233.6 207.4 244.4 ;
      RECT  211.8 254.4 212.6 243.6 ;
      RECT  205.0 254.4 205.8 243.6 ;
      RECT  208.4 244.4 209.2 243.6 ;
      RECT  210.2 254.4 211.0 243.6 ;
      RECT  206.6 254.4 207.4 243.6 ;
      RECT  211.8 254.4 212.6 265.2 ;
      RECT  205.0 254.4 205.8 265.2 ;
      RECT  208.4 264.4 209.2 265.2 ;
      RECT  210.2 254.4 211.0 265.2 ;
      RECT  206.6 254.4 207.4 265.2 ;
      RECT  211.8 275.2 212.6 264.4 ;
      RECT  205.0 275.2 205.8 264.4 ;
      RECT  208.4 265.2 209.2 264.4 ;
      RECT  210.2 275.2 211.0 264.4 ;
      RECT  206.6 275.2 207.4 264.4 ;
      RECT  211.8 275.2 212.6 286.0 ;
      RECT  205.0 275.2 205.8 286.0 ;
      RECT  208.4 285.2 209.2 286.0 ;
      RECT  210.2 275.2 211.0 286.0 ;
      RECT  206.6 275.2 207.4 286.0 ;
      RECT  211.8 296.0 212.6 285.2 ;
      RECT  205.0 296.0 205.8 285.2 ;
      RECT  208.4 286.0 209.2 285.2 ;
      RECT  210.2 296.0 211.0 285.2 ;
      RECT  206.6 296.0 207.4 285.2 ;
      RECT  211.8 296.0 212.6 306.8 ;
      RECT  205.0 296.0 205.8 306.8 ;
      RECT  208.4 306.0 209.2 306.8 ;
      RECT  210.2 296.0 211.0 306.8 ;
      RECT  206.6 296.0 207.4 306.8 ;
      RECT  211.8 316.8 212.6 306.0 ;
      RECT  205.0 316.8 205.8 306.0 ;
      RECT  208.4 306.8 209.2 306.0 ;
      RECT  210.2 316.8 211.0 306.0 ;
      RECT  206.6 316.8 207.4 306.0 ;
      RECT  211.8 316.8 212.6 327.6 ;
      RECT  205.0 316.8 205.8 327.6 ;
      RECT  208.4 326.8 209.2 327.6 ;
      RECT  210.2 316.8 211.0 327.6 ;
      RECT  206.6 316.8 207.4 327.6 ;
      RECT  211.8 337.6 212.6 326.8 ;
      RECT  205.0 337.6 205.8 326.8 ;
      RECT  208.4 327.6 209.2 326.8 ;
      RECT  210.2 337.6 211.0 326.8 ;
      RECT  206.6 337.6 207.4 326.8 ;
      RECT  211.8 337.6 212.6 348.4 ;
      RECT  205.0 337.6 205.8 348.4 ;
      RECT  208.4 347.6 209.2 348.4 ;
      RECT  210.2 337.6 211.0 348.4 ;
      RECT  206.6 337.6 207.4 348.4 ;
      RECT  211.8 358.4 212.6 347.6 ;
      RECT  205.0 358.4 205.8 347.6 ;
      RECT  208.4 348.4 209.2 347.6 ;
      RECT  210.2 358.4 211.0 347.6 ;
      RECT  206.6 358.4 207.4 347.6 ;
      RECT  211.8 358.4 212.6 369.2 ;
      RECT  205.0 358.4 205.8 369.2 ;
      RECT  208.4 368.4 209.2 369.2 ;
      RECT  210.2 358.4 211.0 369.2 ;
      RECT  206.6 358.4 207.4 369.2 ;
      RECT  206.6 171.2 207.4 368.8 ;
      RECT  210.2 171.2 211.0 368.8 ;
      RECT  193.0 171.2 193.8 368.8 ;
      RECT  196.6 171.2 197.4 368.8 ;
      RECT  199.8 171.2 200.6 368.8 ;
      RECT  203.4 171.2 204.2 368.8 ;
      RECT  186.2 171.2 187.0 368.8 ;
      RECT  189.8 171.2 190.6 368.8 ;
      RECT  186.3 154.4 186.9 167.0 ;
      RECT  189.9 154.4 190.5 167.0 ;
      RECT  193.1 154.4 193.7 167.0 ;
      RECT  196.7 154.4 197.3 167.0 ;
      RECT  199.9 154.4 200.5 167.0 ;
      RECT  203.5 154.4 204.1 167.0 ;
      RECT  186.3 154.4 186.9 167.0 ;
      RECT  189.9 154.4 190.5 167.0 ;
      RECT  193.1 154.4 193.7 167.0 ;
      RECT  196.7 154.4 197.3 167.0 ;
      RECT  199.9 154.4 200.5 167.0 ;
      RECT  203.5 154.4 204.1 167.0 ;
      RECT  197.2 130.0 198.0 131.6 ;
      RECT  195.8 126.4 197.0 127.2 ;
      RECT  193.8 126.4 195.2 127.2 ;
      RECT  193.8 127.2 194.6 150.2 ;
      RECT  195.8 127.2 196.6 150.2 ;
      RECT  198.2 143.4 199.0 145.0 ;
      RECT  193.8 117.6 194.6 126.4 ;
      RECT  195.8 117.6 196.6 126.4 ;
      RECT  192.4 117.6 193.2 120.6 ;
      RECT  204.0 130.0 204.8 131.6 ;
      RECT  202.6 126.4 203.8 127.2 ;
      RECT  200.6 126.4 202.0 127.2 ;
      RECT  200.6 127.2 201.4 150.2 ;
      RECT  202.6 127.2 203.4 150.2 ;
      RECT  205.0 143.4 205.8 145.0 ;
      RECT  200.6 117.6 201.4 126.4 ;
      RECT  202.6 117.6 203.4 126.4 ;
      RECT  199.2 117.6 200.0 120.6 ;
      RECT  192.4 117.6 193.2 120.6 ;
      RECT  193.8 127.2 194.6 150.2 ;
      RECT  195.8 127.2 196.6 150.2 ;
      RECT  199.2 117.6 200.0 120.6 ;
      RECT  200.6 127.2 201.4 150.2 ;
      RECT  202.6 127.2 203.4 150.2 ;
      RECT  193.8 111.4 194.6 113.4 ;
      RECT  195.6 85.6 196.4 86.4 ;
      RECT  195.6 79.0 196.4 79.8 ;
      RECT  194.2 104.6 195.0 105.4 ;
      RECT  197.0 90.0 197.8 90.8 ;
      RECT  195.0 96.4 195.8 97.2 ;
      RECT  194.8 72.8 195.6 74.8 ;
      RECT  195.8 108.4 196.6 113.4 ;
      RECT  200.6 111.4 201.4 113.4 ;
      RECT  202.4 85.6 203.2 86.4 ;
      RECT  202.4 79.0 203.2 79.8 ;
      RECT  201.0 104.6 201.8 105.4 ;
      RECT  203.8 90.0 204.6 90.8 ;
      RECT  201.8 96.4 202.6 97.2 ;
      RECT  201.6 72.8 202.4 74.8 ;
      RECT  202.6 108.4 203.4 113.4 ;
      RECT  194.8 72.8 195.6 74.8 ;
      RECT  201.6 72.8 202.4 74.8 ;
      RECT  193.8 111.4 194.6 113.4 ;
      RECT  195.8 108.4 196.6 113.4 ;
      RECT  200.6 111.4 201.4 113.4 ;
      RECT  202.6 108.4 203.4 113.4 ;
      RECT  186.3 167.0 186.9 154.4 ;
      RECT  189.9 167.0 190.5 154.4 ;
      RECT  193.1 167.0 193.7 154.4 ;
      RECT  196.7 167.0 197.3 154.4 ;
      RECT  199.9 167.0 200.5 154.4 ;
      RECT  203.5 167.0 204.1 154.4 ;
      RECT  192.4 120.6 193.2 117.6 ;
      RECT  199.2 120.6 200.0 117.6 ;
      RECT  194.8 74.8 195.6 72.8 ;
      RECT  201.6 74.8 202.4 72.8 ;
      RECT  94.6 193.6 95.2 234.0 ;
      RECT  96.0 193.6 96.6 234.0 ;
      RECT  94.6 235.2 95.2 275.6 ;
      RECT  96.0 235.2 96.6 275.6 ;
      RECT  87.3 192.4 87.9 275.6 ;
      RECT  88.7 192.4 89.3 275.6 ;
      RECT  90.1 192.4 90.7 275.6 ;
      RECT  91.5 192.4 92.1 275.6 ;
      RECT  155.7 192.4 156.3 358.8 ;
      RECT  87.3 192.4 87.9 275.6 ;
      RECT  88.7 192.4 89.3 275.6 ;
      RECT  90.1 192.4 90.7 275.6 ;
      RECT  91.5 192.4 92.1 275.6 ;
      RECT  155.7 192.4 156.3 358.8 ;
      RECT  192.4 117.6 193.2 120.6 ;
      RECT  199.2 117.6 200.0 120.6 ;
      RECT  194.8 72.8 195.6 74.8 ;
      RECT  201.6 72.8 202.4 74.8 ;
      RECT  87.3 192.4 87.9 275.6 ;
      RECT  88.7 192.4 89.3 275.6 ;
      RECT  90.1 192.4 90.7 275.6 ;
      RECT  91.5 192.4 92.1 275.6 ;
      RECT  172.6 72.8 173.2 189.2 ;
      RECT  174.0 72.8 174.6 189.2 ;
      RECT  171.2 72.8 171.8 189.2 ;
      RECT  175.4 72.8 176.0 189.2 ;
      RECT  4.4 3.2 5.2 14.8 ;
      RECT  14.0 3.2 14.8 14.8 ;
      RECT  2.8 6.6 3.6 7.4 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  1.2 5.2 2.0 10.8 ;
      RECT  18.8 9.4 19.6 10.2 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  35.2 7.5 35.8 8.1 ;
      RECT  29.8 10.7 30.4 11.3 ;
      RECT  2.8 6.6 3.6 7.4 ;
      RECT  4.4 36.8 5.2 25.2 ;
      RECT  14.0 36.8 14.8 25.2 ;
      RECT  2.8 33.4 3.6 32.6 ;
      RECT  7.6 31.4 8.4 30.6 ;
      RECT  1.2 34.8 2.0 29.2 ;
      RECT  18.8 30.6 19.6 29.8 ;
      RECT  7.6 31.4 8.4 30.6 ;
      RECT  35.2 32.5 35.8 31.9 ;
      RECT  29.8 29.3 30.4 28.7 ;
      RECT  2.8 33.4 3.6 32.6 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  7.6 30.6 8.4 31.4 ;
      RECT  35.2 7.5 35.8 8.1 ;
      RECT  29.8 10.7 30.4 11.3 ;
      RECT  35.2 31.9 35.8 32.5 ;
      RECT  29.8 28.7 30.4 29.3 ;
      RECT  2.8 0.0 3.4 40.0 ;
      RECT  30.6 162.8 30.0 168.2 ;
      RECT  3.1 162.8 2.5 257.8 ;
      RECT  7.6 8.6 8.4 9.4 ;
      RECT  7.6 30.6 8.4 31.4 ;
      RECT  51.1 0.0 51.7 9.8 ;
      RECT  30.0 162.8 30.6 168.2 ;
      RECT  67.0 293.8 67.8 305.4 ;
      RECT  76.6 293.8 77.4 305.4 ;
      RECT  65.4 297.2 66.2 298.0 ;
      RECT  70.2 299.2 71.0 300.0 ;
      RECT  63.8 295.8 64.6 301.4 ;
      RECT  81.4 300.0 82.2 300.8 ;
      RECT  67.0 327.4 67.8 315.8 ;
      RECT  76.6 327.4 77.4 315.8 ;
      RECT  65.4 324.0 66.2 323.2 ;
      RECT  70.2 322.0 71.0 321.2 ;
      RECT  63.8 325.4 64.6 319.8 ;
      RECT  81.4 321.2 82.2 320.4 ;
      RECT  67.0 333.8 67.8 345.4 ;
      RECT  76.6 333.8 77.4 345.4 ;
      RECT  65.4 337.2 66.2 338.0 ;
      RECT  70.2 339.2 71.0 340.0 ;
      RECT  63.8 335.8 64.6 341.4 ;
      RECT  81.4 340.0 82.2 340.8 ;
      RECT  67.0 367.4 67.8 355.8 ;
      RECT  76.6 367.4 77.4 355.8 ;
      RECT  65.4 364.0 66.2 363.2 ;
      RECT  70.2 362.0 71.0 361.2 ;
      RECT  63.8 365.4 64.6 359.8 ;
      RECT  81.4 361.2 82.2 360.4 ;
      RECT  70.2 299.2 71.0 300.0 ;
      RECT  70.2 321.2 71.0 322.0 ;
      RECT  70.2 339.2 71.0 340.0 ;
      RECT  70.2 361.2 71.0 362.0 ;
      RECT  81.4 300.0 82.2 300.8 ;
      RECT  81.4 320.4 82.2 321.2 ;
      RECT  81.4 340.0 82.2 340.8 ;
      RECT  81.4 360.4 82.2 361.2 ;
      RECT  182.6 49.0 183.4 60.6 ;
      RECT  192.2 49.0 193.0 60.6 ;
      RECT  181.0 52.4 181.8 53.2 ;
      RECT  185.8 54.4 186.6 55.2 ;
      RECT  179.4 51.0 180.2 56.6 ;
      RECT  197.0 55.2 197.8 56.0 ;
      RECT  204.4 49.0 205.2 60.6 ;
      RECT  214.0 49.0 214.8 60.6 ;
      RECT  202.8 52.4 203.6 53.2 ;
      RECT  207.6 54.4 208.4 55.2 ;
      RECT  201.2 51.0 202.0 56.6 ;
      RECT  218.8 55.2 219.6 56.0 ;
      RECT  185.8 54.4 186.6 55.2 ;
      RECT  207.6 54.4 208.4 55.2 ;
      RECT  197.0 55.2 197.8 56.0 ;
      RECT  218.8 55.2 219.6 56.0 ;
   LAYER  m3 ;
      RECT  194.8 222.8 195.6 223.6 ;
      RECT  194.8 202.0 195.6 202.8 ;
      RECT  201.6 243.6 202.4 244.4 ;
      RECT  201.6 243.6 202.4 244.4 ;
      RECT  201.6 264.4 202.4 265.2 ;
      RECT  201.6 285.2 202.4 286.0 ;
      RECT  201.6 202.0 202.4 202.8 ;
      RECT  201.6 326.8 202.4 327.6 ;
      RECT  201.6 326.8 202.4 327.6 ;
      RECT  201.6 347.6 202.4 348.4 ;
      RECT  194.8 347.6 195.6 348.4 ;
      RECT  194.8 243.6 195.6 244.4 ;
      RECT  194.8 243.6 195.6 244.4 ;
      RECT  201.6 306.0 202.4 306.8 ;
      RECT  194.8 326.8 195.6 327.6 ;
      RECT  194.8 306.0 195.6 306.8 ;
      RECT  194.8 264.4 195.6 265.2 ;
      RECT  194.8 326.8 195.6 327.6 ;
      RECT  194.8 285.2 195.6 286.0 ;
      RECT  201.6 222.8 202.4 223.6 ;
      RECT  205.0 197.0 205.8 197.8 ;
      RECT  198.2 238.6 199.0 239.4 ;
      RECT  191.4 207.0 192.2 207.8 ;
      RECT  198.2 352.6 199.0 353.4 ;
      RECT  198.2 342.6 199.0 343.4 ;
      RECT  191.4 290.2 192.2 291.0 ;
      RECT  191.4 259.4 192.2 260.2 ;
      RECT  198.2 301.0 199.0 301.8 ;
      RECT  198.2 331.8 199.0 332.6 ;
      RECT  205.0 352.6 205.8 353.4 ;
      RECT  205.0 301.0 205.8 301.8 ;
      RECT  191.4 311.0 192.2 311.8 ;
      RECT  198.2 269.4 199.0 270.2 ;
      RECT  198.2 207.0 199.0 207.8 ;
      RECT  205.0 290.2 205.8 291.0 ;
      RECT  191.4 301.0 192.2 301.8 ;
      RECT  205.0 269.4 205.8 270.2 ;
      RECT  205.0 238.6 205.8 239.4 ;
      RECT  198.2 227.8 199.0 228.6 ;
      RECT  191.4 227.8 192.2 228.6 ;
      RECT  191.4 197.0 192.2 197.8 ;
      RECT  191.4 248.6 192.2 249.4 ;
      RECT  198.2 248.6 199.0 249.4 ;
      RECT  191.4 321.8 192.2 322.6 ;
      RECT  205.0 321.8 205.8 322.6 ;
      RECT  198.2 217.8 199.0 218.6 ;
      RECT  198.2 290.2 199.0 291.0 ;
      RECT  191.4 342.6 192.2 343.4 ;
      RECT  205.0 248.6 205.8 249.4 ;
      RECT  205.0 311.0 205.8 311.8 ;
      RECT  191.4 352.6 192.2 353.4 ;
      RECT  191.4 217.8 192.2 218.6 ;
      RECT  205.0 280.2 205.8 281.0 ;
      RECT  205.0 207.0 205.8 207.8 ;
      RECT  205.0 217.8 205.8 218.6 ;
      RECT  198.2 321.8 199.0 322.6 ;
      RECT  205.0 259.4 205.8 260.2 ;
      RECT  191.4 238.6 192.2 239.4 ;
      RECT  198.2 280.2 199.0 281.0 ;
      RECT  191.4 331.8 192.2 332.6 ;
      RECT  191.4 269.4 192.2 270.2 ;
      RECT  191.4 280.2 192.2 281.0 ;
      RECT  205.0 342.6 205.8 343.4 ;
      RECT  198.2 197.0 199.0 197.8 ;
      RECT  205.0 331.8 205.8 332.6 ;
      RECT  198.2 259.4 199.0 260.2 ;
      RECT  205.0 227.8 205.8 228.6 ;
      RECT  198.2 311.0 199.0 311.8 ;
      RECT  194.8 182.0 195.6 181.2 ;
      RECT  201.6 182.0 202.4 181.2 ;
      RECT  198.2 187.0 199.0 186.2 ;
      RECT  191.4 187.0 192.2 186.2 ;
      RECT  205.0 187.0 205.8 186.2 ;
      RECT  194.8 181.2 195.6 182.0 ;
      RECT  201.6 181.2 202.4 182.0 ;
      RECT  198.2 176.2 199.0 177.0 ;
      RECT  191.4 176.2 192.2 177.0 ;
      RECT  205.0 176.2 205.8 177.0 ;
      RECT  194.8 368.4 195.6 369.2 ;
      RECT  201.6 368.4 202.4 369.2 ;
      RECT  198.2 363.4 199.0 364.2 ;
      RECT  191.4 363.4 192.2 364.2 ;
      RECT  205.0 363.4 205.8 364.2 ;
      RECT  181.2 347.6 182.0 348.4 ;
      RECT  181.2 222.8 182.0 223.6 ;
      RECT  181.2 202.0 182.0 202.8 ;
      RECT  181.2 222.8 182.0 223.6 ;
      RECT  181.2 368.4 182.0 369.2 ;
      RECT  181.2 181.2 182.0 182.0 ;
      RECT  181.2 306.0 182.0 306.8 ;
      RECT  181.2 285.2 182.0 286.0 ;
      RECT  181.2 243.6 182.0 244.4 ;
      RECT  181.2 306.0 182.0 306.8 ;
      RECT  181.2 264.4 182.0 265.2 ;
      RECT  181.2 326.8 182.0 327.6 ;
      RECT  184.6 217.8 185.4 218.6 ;
      RECT  184.6 331.8 185.4 332.6 ;
      RECT  177.8 186.2 178.6 187.0 ;
      RECT  184.6 363.4 185.4 364.2 ;
      RECT  184.6 321.8 185.4 322.6 ;
      RECT  177.8 269.4 178.6 270.2 ;
      RECT  177.8 238.6 178.6 239.4 ;
      RECT  184.6 280.2 185.4 281.0 ;
      RECT  184.6 311.0 185.4 311.8 ;
      RECT  184.6 342.6 185.4 343.4 ;
      RECT  177.8 290.2 178.6 291.0 ;
      RECT  184.6 248.6 185.4 249.4 ;
      RECT  184.6 186.2 185.4 187.0 ;
      RECT  177.8 280.2 178.6 281.0 ;
      RECT  184.6 207.0 185.4 207.8 ;
      RECT  177.8 176.2 178.6 177.0 ;
      RECT  177.8 207.0 178.6 207.8 ;
      RECT  177.8 227.8 178.6 228.6 ;
      RECT  184.6 227.8 185.4 228.6 ;
      RECT  177.8 301.0 178.6 301.8 ;
      RECT  184.6 197.0 185.4 197.8 ;
      RECT  184.6 269.4 185.4 270.2 ;
      RECT  177.8 321.8 178.6 322.6 ;
      RECT  177.8 331.8 178.6 332.6 ;
      RECT  177.8 197.0 178.6 197.8 ;
      RECT  184.6 352.6 185.4 353.4 ;
      RECT  177.8 363.4 178.6 364.2 ;
      RECT  184.6 301.0 185.4 301.8 ;
      RECT  177.8 217.8 178.6 218.6 ;
      RECT  177.8 352.6 178.6 353.4 ;
      RECT  184.6 259.4 185.4 260.2 ;
      RECT  177.8 311.0 178.6 311.8 ;
      RECT  177.8 248.6 178.6 249.4 ;
      RECT  177.8 259.4 178.6 260.2 ;
      RECT  177.8 342.6 178.6 343.4 ;
      RECT  184.6 176.2 185.4 177.0 ;
      RECT  184.6 238.6 185.4 239.4 ;
      RECT  184.6 290.2 185.4 291.0 ;
      RECT  208.4 347.6 209.2 348.4 ;
      RECT  208.4 222.8 209.2 223.6 ;
      RECT  208.4 202.0 209.2 202.8 ;
      RECT  208.4 222.8 209.2 223.6 ;
      RECT  208.4 368.4 209.2 369.2 ;
      RECT  208.4 181.2 209.2 182.0 ;
      RECT  208.4 306.0 209.2 306.8 ;
      RECT  208.4 285.2 209.2 286.0 ;
      RECT  208.4 243.6 209.2 244.4 ;
      RECT  208.4 306.0 209.2 306.8 ;
      RECT  208.4 264.4 209.2 265.2 ;
      RECT  208.4 326.8 209.2 327.6 ;
      RECT  211.8 217.8 212.6 218.6 ;
      RECT  211.8 331.8 212.6 332.6 ;
      RECT  205.0 186.2 205.8 187.0 ;
      RECT  211.8 363.4 212.6 364.2 ;
      RECT  211.8 321.8 212.6 322.6 ;
      RECT  205.0 269.4 205.8 270.2 ;
      RECT  205.0 238.6 205.8 239.4 ;
      RECT  211.8 280.2 212.6 281.0 ;
      RECT  211.8 311.0 212.6 311.8 ;
      RECT  211.8 342.6 212.6 343.4 ;
      RECT  205.0 290.2 205.8 291.0 ;
      RECT  211.8 248.6 212.6 249.4 ;
      RECT  211.8 186.2 212.6 187.0 ;
      RECT  205.0 280.2 205.8 281.0 ;
      RECT  211.8 207.0 212.6 207.8 ;
      RECT  205.0 176.2 205.8 177.0 ;
      RECT  205.0 207.0 205.8 207.8 ;
      RECT  205.0 227.8 205.8 228.6 ;
      RECT  211.8 227.8 212.6 228.6 ;
      RECT  205.0 301.0 205.8 301.8 ;
      RECT  211.8 197.0 212.6 197.8 ;
      RECT  211.8 269.4 212.6 270.2 ;
      RECT  205.0 321.8 205.8 322.6 ;
      RECT  205.0 331.8 205.8 332.6 ;
      RECT  205.0 197.0 205.8 197.8 ;
      RECT  211.8 352.6 212.6 353.4 ;
      RECT  205.0 363.4 205.8 364.2 ;
      RECT  211.8 301.0 212.6 301.8 ;
      RECT  205.0 217.8 205.8 218.6 ;
      RECT  205.0 352.6 205.8 353.4 ;
      RECT  211.8 259.4 212.6 260.2 ;
      RECT  205.0 311.0 205.8 311.8 ;
      RECT  205.0 248.6 205.8 249.4 ;
      RECT  205.0 259.4 205.8 260.2 ;
      RECT  205.0 342.6 205.8 343.4 ;
      RECT  211.8 176.2 212.6 177.0 ;
      RECT  211.8 238.6 212.6 239.4 ;
      RECT  211.8 290.2 212.6 291.0 ;
      RECT  181.3 285.3 181.9 285.9 ;
      RECT  194.9 202.1 195.5 202.7 ;
      RECT  188.0 222.8 188.8 223.6 ;
      RECT  208.5 347.7 209.1 348.3 ;
      RECT  208.5 181.3 209.1 181.9 ;
      RECT  194.9 306.1 195.5 306.7 ;
      RECT  188.0 243.6 188.8 244.4 ;
      RECT  201.7 368.5 202.3 369.1 ;
      RECT  181.3 368.5 181.9 369.1 ;
      RECT  194.9 326.9 195.5 327.5 ;
      RECT  201.7 202.1 202.3 202.7 ;
      RECT  208.5 222.9 209.1 223.5 ;
      RECT  181.3 202.1 181.9 202.7 ;
      RECT  188.0 347.6 188.8 348.4 ;
      RECT  188.0 264.4 188.8 265.2 ;
      RECT  194.9 264.5 195.5 265.1 ;
      RECT  201.7 285.3 202.3 285.9 ;
      RECT  181.3 306.1 181.9 306.7 ;
      RECT  201.7 243.7 202.3 244.3 ;
      RECT  194.9 285.3 195.5 285.9 ;
      RECT  194.9 222.9 195.5 223.5 ;
      RECT  188.0 181.2 188.8 182.0 ;
      RECT  188.0 306.0 188.8 306.8 ;
      RECT  201.7 347.7 202.3 348.3 ;
      RECT  188.0 326.8 188.8 327.6 ;
      RECT  208.5 285.3 209.1 285.9 ;
      RECT  181.3 222.9 181.9 223.5 ;
      RECT  194.9 347.7 195.5 348.3 ;
      RECT  181.3 326.9 181.9 327.5 ;
      RECT  201.7 222.9 202.3 223.5 ;
      RECT  201.7 264.5 202.3 265.1 ;
      RECT  181.3 181.3 181.9 181.9 ;
      RECT  208.5 368.5 209.1 369.1 ;
      RECT  208.5 306.1 209.1 306.7 ;
      RECT  208.5 326.9 209.1 327.5 ;
      RECT  181.3 347.7 181.9 348.3 ;
      RECT  194.9 243.7 195.5 244.3 ;
      RECT  201.7 326.9 202.3 327.5 ;
      RECT  194.9 368.5 195.5 369.1 ;
      RECT  188.0 285.2 188.8 286.0 ;
      RECT  208.5 202.1 209.1 202.7 ;
      RECT  208.5 264.5 209.1 265.1 ;
      RECT  201.7 306.1 202.3 306.7 ;
      RECT  194.9 181.3 195.5 181.9 ;
      RECT  181.3 243.7 181.9 244.3 ;
      RECT  188.0 368.4 188.8 369.2 ;
      RECT  181.3 264.5 181.9 265.1 ;
      RECT  188.0 202.0 188.8 202.8 ;
      RECT  208.5 243.7 209.1 244.3 ;
      RECT  201.7 181.3 202.3 181.9 ;
      RECT  184.6 217.8 185.4 218.6 ;
      RECT  191.5 280.3 192.1 280.9 ;
      RECT  191.4 280.2 192.2 281.0 ;
      RECT  177.9 311.1 178.5 311.7 ;
      RECT  205.1 290.3 205.7 290.9 ;
      RECT  198.3 238.7 198.9 239.3 ;
      RECT  211.9 321.9 212.5 322.5 ;
      RECT  191.4 352.6 192.2 353.4 ;
      RECT  177.9 259.5 178.5 260.1 ;
      RECT  205.1 280.3 205.7 280.9 ;
      RECT  191.4 342.6 192.2 343.4 ;
      RECT  191.5 363.5 192.1 364.1 ;
      RECT  211.9 352.7 212.5 353.3 ;
      RECT  198.3 207.1 198.9 207.7 ;
      RECT  184.7 331.9 185.3 332.5 ;
      RECT  191.4 301.0 192.2 301.8 ;
      RECT  184.7 311.1 185.3 311.7 ;
      RECT  198.3 311.1 198.9 311.7 ;
      RECT  184.7 186.3 185.3 186.9 ;
      RECT  184.7 176.3 185.3 176.9 ;
      RECT  211.9 301.1 212.5 301.7 ;
      RECT  198.3 363.5 198.9 364.1 ;
      RECT  184.7 207.1 185.3 207.7 ;
      RECT  191.4 290.2 192.2 291.0 ;
      RECT  205.1 352.7 205.7 353.3 ;
      RECT  198.3 259.5 198.9 260.1 ;
      RECT  191.5 269.5 192.1 270.1 ;
      RECT  191.5 197.1 192.1 197.7 ;
      RECT  211.9 238.7 212.5 239.3 ;
      RECT  184.7 363.5 185.3 364.1 ;
      RECT  177.9 301.1 178.5 301.7 ;
      RECT  198.3 217.9 198.9 218.5 ;
      RECT  205.1 197.1 205.7 197.7 ;
      RECT  177.9 176.3 178.5 176.9 ;
      RECT  211.9 290.3 212.5 290.9 ;
      RECT  177.9 238.7 178.5 239.3 ;
      RECT  184.6 176.2 185.4 177.0 ;
      RECT  198.3 227.9 198.9 228.5 ;
      RECT  184.7 290.3 185.3 290.9 ;
      RECT  191.5 248.7 192.1 249.3 ;
      RECT  211.9 197.1 212.5 197.7 ;
      RECT  191.5 301.1 192.1 301.7 ;
      RECT  205.1 238.7 205.7 239.3 ;
      RECT  205.1 248.7 205.7 249.3 ;
      RECT  198.3 301.1 198.9 301.7 ;
      RECT  184.6 342.6 185.4 343.4 ;
      RECT  205.1 259.5 205.7 260.1 ;
      RECT  191.5 176.3 192.1 176.9 ;
      RECT  211.9 363.5 212.5 364.1 ;
      RECT  205.1 186.3 205.7 186.9 ;
      RECT  184.6 186.2 185.4 187.0 ;
      RECT  211.9 186.3 212.5 186.9 ;
      RECT  191.4 269.4 192.2 270.2 ;
      RECT  198.3 352.7 198.9 353.3 ;
      RECT  205.1 301.1 205.7 301.7 ;
      RECT  191.5 321.9 192.1 322.5 ;
      RECT  205.1 301.1 205.7 301.7 ;
      RECT  184.7 342.7 185.3 343.3 ;
      RECT  184.6 207.0 185.4 207.8 ;
      RECT  191.5 227.9 192.1 228.5 ;
      RECT  184.6 227.8 185.4 228.6 ;
      RECT  205.1 311.1 205.7 311.7 ;
      RECT  184.7 352.7 185.3 353.3 ;
      RECT  205.1 311.1 205.7 311.7 ;
      RECT  211.9 217.9 212.5 218.5 ;
      RECT  191.5 217.9 192.1 218.5 ;
      RECT  191.4 227.8 192.2 228.6 ;
      RECT  198.3 197.1 198.9 197.7 ;
      RECT  191.4 197.0 192.2 197.8 ;
      RECT  184.7 321.9 185.3 322.5 ;
      RECT  177.9 248.7 178.5 249.3 ;
      RECT  177.9 352.7 178.5 353.3 ;
      RECT  205.1 269.5 205.7 270.1 ;
      RECT  177.9 342.7 178.5 343.3 ;
      RECT  191.5 331.9 192.1 332.5 ;
      RECT  198.3 331.9 198.9 332.5 ;
      RECT  191.4 321.8 192.2 322.6 ;
      RECT  184.6 238.6 185.4 239.4 ;
      RECT  184.6 290.2 185.4 291.0 ;
      RECT  184.7 280.3 185.3 280.9 ;
      RECT  205.1 331.9 205.7 332.5 ;
      RECT  191.4 176.2 192.2 177.0 ;
      RECT  184.7 259.5 185.3 260.1 ;
      RECT  211.9 280.3 212.5 280.9 ;
      RECT  198.3 290.3 198.9 290.9 ;
      RECT  184.6 321.8 185.4 322.6 ;
      RECT  177.9 280.3 178.5 280.9 ;
      RECT  211.9 342.7 212.5 343.3 ;
      RECT  211.9 227.9 212.5 228.5 ;
      RECT  184.6 280.2 185.4 281.0 ;
      RECT  184.7 197.1 185.3 197.7 ;
      RECT  198.3 248.7 198.9 249.3 ;
      RECT  184.7 248.7 185.3 249.3 ;
      RECT  184.6 248.6 185.4 249.4 ;
      RECT  205.1 176.3 205.7 176.9 ;
      RECT  177.9 321.9 178.5 322.5 ;
      RECT  198.3 342.7 198.9 343.3 ;
      RECT  205.1 227.9 205.7 228.5 ;
      RECT  205.1 227.9 205.7 228.5 ;
      RECT  191.4 217.8 192.2 218.6 ;
      RECT  211.9 176.3 212.5 176.9 ;
      RECT  184.6 269.4 185.4 270.2 ;
      RECT  184.7 227.9 185.3 228.5 ;
      RECT  191.5 290.3 192.1 290.9 ;
      RECT  198.3 186.3 198.9 186.9 ;
      RECT  191.5 311.1 192.1 311.7 ;
      RECT  198.3 269.5 198.9 270.1 ;
      RECT  184.6 301.0 185.4 301.8 ;
      RECT  211.9 269.5 212.5 270.1 ;
      RECT  191.4 238.6 192.2 239.4 ;
      RECT  205.1 207.1 205.7 207.7 ;
      RECT  191.5 238.7 192.1 239.3 ;
      RECT  191.4 363.4 192.2 364.2 ;
      RECT  177.9 227.9 178.5 228.5 ;
      RECT  177.9 197.1 178.5 197.7 ;
      RECT  211.9 248.7 212.5 249.3 ;
      RECT  191.4 311.0 192.2 311.8 ;
      RECT  177.9 331.9 178.5 332.5 ;
      RECT  184.7 301.1 185.3 301.7 ;
      RECT  184.6 363.4 185.4 364.2 ;
      RECT  184.6 331.8 185.4 332.6 ;
      RECT  184.6 311.0 185.4 311.8 ;
      RECT  177.9 290.3 178.5 290.9 ;
      RECT  205.1 321.9 205.7 322.5 ;
      RECT  211.9 207.1 212.5 207.7 ;
      RECT  184.7 217.9 185.3 218.5 ;
      RECT  205.1 217.9 205.7 218.5 ;
      RECT  191.4 248.6 192.2 249.4 ;
      RECT  177.9 217.9 178.5 218.5 ;
      RECT  191.5 207.1 192.1 207.7 ;
      RECT  211.9 259.5 212.5 260.1 ;
      RECT  198.3 280.3 198.9 280.9 ;
      RECT  184.6 197.0 185.4 197.8 ;
      RECT  177.9 269.5 178.5 270.1 ;
      RECT  205.1 363.5 205.7 364.1 ;
      RECT  191.5 259.5 192.1 260.1 ;
      RECT  211.9 311.1 212.5 311.7 ;
      RECT  198.3 321.9 198.9 322.5 ;
      RECT  184.7 269.5 185.3 270.1 ;
      RECT  205.1 342.7 205.7 343.3 ;
      RECT  191.4 259.4 192.2 260.2 ;
      RECT  191.4 186.2 192.2 187.0 ;
      RECT  184.7 238.7 185.3 239.3 ;
      RECT  184.6 259.4 185.4 260.2 ;
      RECT  177.9 363.5 178.5 364.1 ;
      RECT  191.5 186.3 192.1 186.9 ;
      RECT  191.5 342.7 192.1 343.3 ;
      RECT  191.5 352.7 192.1 353.3 ;
      RECT  198.3 176.3 198.9 176.9 ;
      RECT  177.9 186.3 178.5 186.9 ;
      RECT  211.9 331.9 212.5 332.5 ;
      RECT  191.4 331.8 192.2 332.6 ;
      RECT  177.9 207.1 178.5 207.7 ;
      RECT  184.6 352.6 185.4 353.4 ;
      RECT  191.4 207.0 192.2 207.8 ;
      RECT  187.8 160.8 188.6 161.6 ;
      RECT  194.6 160.8 195.4 161.6 ;
      RECT  201.4 160.8 202.2 161.6 ;
      RECT  201.4 160.8 202.2 161.6 ;
      RECT  194.6 160.8 195.4 161.6 ;
      RECT  187.8 160.8 188.6 161.6 ;
      RECT  204.0 130.4 204.8 131.2 ;
      RECT  197.2 130.4 198.0 131.2 ;
      RECT  205.0 143.8 205.8 144.6 ;
      RECT  198.2 143.8 199.0 144.6 ;
      RECT  201.8 96.4 202.6 97.2 ;
      RECT  195.0 96.4 195.8 97.2 ;
      RECT  195.6 79.0 196.4 79.8 ;
      RECT  202.4 79.0 203.2 79.8 ;
      RECT  201.0 104.6 201.8 105.4 ;
      RECT  195.6 85.6 196.4 86.4 ;
      RECT  202.4 85.6 203.2 86.4 ;
      RECT  197.0 90.0 197.8 90.8 ;
      RECT  203.8 90.0 204.6 90.8 ;
      RECT  194.2 104.6 195.0 105.4 ;
      RECT  187.8 161.6 188.6 160.8 ;
      RECT  197.2 131.2 198.0 130.4 ;
      RECT  194.6 161.6 195.4 160.8 ;
      RECT  204.0 131.2 204.8 130.4 ;
      RECT  202.4 79.8 203.2 79.0 ;
      RECT  201.8 97.2 202.6 96.4 ;
      RECT  195.6 79.8 196.4 79.0 ;
      RECT  201.4 161.6 202.2 160.8 ;
      RECT  195.0 97.2 195.8 96.4 ;
      RECT  198.2 144.6 199.0 143.8 ;
      RECT  202.4 86.4 203.2 85.6 ;
      RECT  201.0 105.4 201.8 104.6 ;
      RECT  194.2 105.4 195.0 104.6 ;
      RECT  205.0 144.6 205.8 143.8 ;
      RECT  197.0 90.8 197.8 90.0 ;
      RECT  203.8 90.8 204.6 90.0 ;
      RECT  195.6 86.4 196.4 85.6 ;
      RECT  118.7 223.2 119.5 224.0 ;
      RECT  118.7 223.2 119.5 224.0 ;
      RECT  103.7 223.2 104.5 224.0 ;
      RECT  103.7 223.2 104.5 224.0 ;
      RECT  118.7 202.4 119.5 203.2 ;
      RECT  118.7 202.4 119.5 203.2 ;
      RECT  103.7 202.4 104.5 203.2 ;
      RECT  103.7 202.4 104.5 203.2 ;
      RECT  103.7 192.0 104.5 192.8 ;
      RECT  118.7 233.6 119.5 234.4 ;
      RECT  118.7 192.0 119.5 192.8 ;
      RECT  118.7 212.8 119.5 213.6 ;
      RECT  103.7 233.6 104.5 234.4 ;
      RECT  103.7 212.8 104.5 213.6 ;
      RECT  118.7 264.8 119.5 265.6 ;
      RECT  118.7 264.8 119.5 265.6 ;
      RECT  103.7 264.8 104.5 265.6 ;
      RECT  103.7 264.8 104.5 265.6 ;
      RECT  118.7 244.0 119.5 244.8 ;
      RECT  118.7 244.0 119.5 244.8 ;
      RECT  103.7 244.0 104.5 244.8 ;
      RECT  103.7 244.0 104.5 244.8 ;
      RECT  103.7 233.6 104.5 234.4 ;
      RECT  118.7 275.2 119.5 276.0 ;
      RECT  118.7 233.6 119.5 234.4 ;
      RECT  118.7 254.4 119.5 255.2 ;
      RECT  103.7 275.2 104.5 276.0 ;
      RECT  103.7 254.4 104.5 255.2 ;
      RECT  144.7 244.0 145.5 244.8 ;
      RECT  144.7 264.8 145.5 265.6 ;
      RECT  144.7 264.8 145.5 265.6 ;
      RECT  144.7 202.4 145.5 203.2 ;
      RECT  144.7 202.4 145.5 203.2 ;
      RECT  118.7 264.8 119.5 265.6 ;
      RECT  144.7 348.0 145.5 348.8 ;
      RECT  103.7 244.0 104.5 244.8 ;
      RECT  118.7 244.0 119.5 244.8 ;
      RECT  144.7 223.2 145.5 224.0 ;
      RECT  144.7 223.2 145.5 224.0 ;
      RECT  118.7 202.4 119.5 203.2 ;
      RECT  144.7 327.2 145.5 328.0 ;
      RECT  103.7 264.8 104.5 265.6 ;
      RECT  103.7 202.4 104.5 203.2 ;
      RECT  103.7 223.2 104.5 224.0 ;
      RECT  118.7 223.2 119.5 224.0 ;
      RECT  144.7 306.4 145.5 307.2 ;
      RECT  144.7 285.6 145.5 286.4 ;
      RECT  144.7 285.6 145.5 286.4 ;
      RECT  103.7 254.4 104.5 255.2 ;
      RECT  144.7 296.0 145.5 296.8 ;
      RECT  118.7 254.4 119.5 255.2 ;
      RECT  118.7 233.6 119.5 234.4 ;
      RECT  144.7 358.4 145.5 359.2 ;
      RECT  144.7 192.0 145.5 192.8 ;
      RECT  144.7 212.8 145.5 213.6 ;
      RECT  144.7 337.6 145.5 338.4 ;
      RECT  103.7 192.0 104.5 192.8 ;
      RECT  118.7 192.0 119.5 192.8 ;
      RECT  144.7 275.2 145.5 276.0 ;
      RECT  144.7 316.8 145.5 317.6 ;
      RECT  144.7 254.4 145.5 255.2 ;
      RECT  118.7 212.8 119.5 213.6 ;
      RECT  103.7 233.6 104.5 234.4 ;
      RECT  103.7 275.2 104.5 276.0 ;
      RECT  103.7 212.8 104.5 213.6 ;
      RECT  118.7 275.2 119.5 276.0 ;
      RECT  144.7 233.6 145.5 234.4 ;
      RECT  165.5 223.2 166.3 224.0 ;
      RECT  165.5 306.4 166.3 307.2 ;
      RECT  165.5 348.0 166.3 348.8 ;
      RECT  165.5 244.0 166.3 244.8 ;
      RECT  165.5 202.4 166.3 203.2 ;
      RECT  165.5 285.6 166.3 286.4 ;
      RECT  165.5 285.6 166.3 286.4 ;
      RECT  165.5 264.8 166.3 265.6 ;
      RECT  165.5 327.2 166.3 328.0 ;
      RECT  165.5 202.4 166.3 203.2 ;
      RECT  165.5 223.2 166.3 224.0 ;
      RECT  165.5 264.8 166.3 265.6 ;
      RECT  165.5 358.4 166.3 359.2 ;
      RECT  165.5 254.4 166.3 255.2 ;
      RECT  165.5 275.2 166.3 276.0 ;
      RECT  165.5 296.0 166.3 296.8 ;
      RECT  165.5 316.8 166.3 317.6 ;
      RECT  165.5 192.0 166.3 192.8 ;
      RECT  165.5 233.6 166.3 234.4 ;
      RECT  165.5 212.8 166.3 213.6 ;
      RECT  165.5 337.6 166.3 338.4 ;
      RECT  103.7 244.0 104.5 244.8 ;
      RECT  165.5 348.0 166.3 348.8 ;
      RECT  165.5 264.8 166.3 265.6 ;
      RECT  144.7 202.4 145.5 203.2 ;
      RECT  165.5 223.2 166.3 224.0 ;
      RECT  118.7 264.8 119.5 265.6 ;
      RECT  144.7 327.2 145.5 328.0 ;
      RECT  118.7 244.0 119.5 244.8 ;
      RECT  165.5 327.2 166.3 328.0 ;
      RECT  144.7 348.0 145.5 348.8 ;
      RECT  118.7 202.4 119.5 203.2 ;
      RECT  103.7 264.8 104.5 265.6 ;
      RECT  165.5 285.6 166.3 286.4 ;
      RECT  165.5 202.4 166.3 203.2 ;
      RECT  103.7 223.2 104.5 224.0 ;
      RECT  144.7 223.2 145.5 224.0 ;
      RECT  144.7 244.0 145.5 244.8 ;
      RECT  165.5 244.0 166.3 244.8 ;
      RECT  144.7 306.4 145.5 307.2 ;
      RECT  118.7 223.2 119.5 224.0 ;
      RECT  103.7 202.4 104.5 203.2 ;
      RECT  165.5 306.4 166.3 307.2 ;
      RECT  144.7 264.8 145.5 265.6 ;
      RECT  144.7 285.6 145.5 286.4 ;
      RECT  165.5 192.0 166.3 192.8 ;
      RECT  118.7 192.0 119.5 192.8 ;
      RECT  103.7 254.4 104.5 255.2 ;
      RECT  103.7 233.6 104.5 234.4 ;
      RECT  118.7 275.2 119.5 276.0 ;
      RECT  165.5 337.6 166.3 338.4 ;
      RECT  144.7 254.4 145.5 255.2 ;
      RECT  165.5 275.2 166.3 276.0 ;
      RECT  165.5 358.4 166.3 359.2 ;
      RECT  144.7 296.0 145.5 296.8 ;
      RECT  144.7 358.4 145.5 359.2 ;
      RECT  165.5 212.8 166.3 213.6 ;
      RECT  144.7 233.6 145.5 234.4 ;
      RECT  165.5 254.4 166.3 255.2 ;
      RECT  103.7 192.0 104.5 192.8 ;
      RECT  144.7 192.0 145.5 192.8 ;
      RECT  144.7 275.2 145.5 276.0 ;
      RECT  103.7 275.2 104.5 276.0 ;
      RECT  118.7 233.6 119.5 234.4 ;
      RECT  144.7 316.8 145.5 317.6 ;
      RECT  165.5 296.0 166.3 296.8 ;
      RECT  144.7 337.6 145.5 338.4 ;
      RECT  165.5 233.6 166.3 234.4 ;
      RECT  144.7 212.8 145.5 213.6 ;
      RECT  165.5 316.8 166.3 317.6 ;
      RECT  118.7 212.8 119.5 213.6 ;
      RECT  118.7 254.4 119.5 255.2 ;
      RECT  103.7 212.8 104.5 213.6 ;
      RECT  165.5 202.4 166.3 203.2 ;
      RECT  103.7 223.2 104.5 224.0 ;
      RECT  188.0 222.8 188.8 223.6 ;
      RECT  118.7 264.8 119.5 265.6 ;
      RECT  208.5 181.3 209.1 181.9 ;
      RECT  194.9 326.9 195.5 327.5 ;
      RECT  103.7 264.8 104.5 265.6 ;
      RECT  144.7 348.0 145.5 348.8 ;
      RECT  181.3 306.1 181.9 306.7 ;
      RECT  201.7 243.7 202.3 244.3 ;
      RECT  194.9 285.3 195.5 285.9 ;
      RECT  194.9 347.7 195.5 348.3 ;
      RECT  208.5 306.1 209.1 306.7 ;
      RECT  195.0 96.4 195.8 97.2 ;
      RECT  144.7 202.4 145.5 203.2 ;
      RECT  201.8 96.4 202.6 97.2 ;
      RECT  165.5 244.0 166.3 244.8 ;
      RECT  103.7 244.0 104.5 244.8 ;
      RECT  187.8 160.8 188.6 161.6 ;
      RECT  144.7 306.4 145.5 307.2 ;
      RECT  188.0 243.6 188.8 244.4 ;
      RECT  188.0 347.6 188.8 348.4 ;
      RECT  188.0 264.4 188.8 265.2 ;
      RECT  201.7 285.3 202.3 285.9 ;
      RECT  194.9 222.9 195.5 223.5 ;
      RECT  188.0 326.8 188.8 327.6 ;
      RECT  181.3 222.9 181.9 223.5 ;
      RECT  181.3 326.9 181.9 327.5 ;
      RECT  194.9 368.5 195.5 369.1 ;
      RECT  144.7 223.2 145.5 224.0 ;
      RECT  201.7 306.1 202.3 306.7 ;
      RECT  194.9 181.3 195.5 181.9 ;
      RECT  188.0 202.0 188.8 202.8 ;
      RECT  208.5 243.7 209.1 244.3 ;
      RECT  181.3 368.5 181.9 369.1 ;
      RECT  201.7 181.3 202.3 181.9 ;
      RECT  165.5 306.4 166.3 307.2 ;
      RECT  165.5 223.2 166.3 224.0 ;
      RECT  181.3 285.3 181.9 285.9 ;
      RECT  201.7 368.5 202.3 369.1 ;
      RECT  194.9 306.1 195.5 306.7 ;
      RECT  165.5 285.6 166.3 286.4 ;
      RECT  208.5 222.9 209.1 223.5 ;
      RECT  194.9 264.5 195.5 265.1 ;
      RECT  188.0 181.2 188.8 182.0 ;
      RECT  201.7 347.7 202.3 348.3 ;
      RECT  208.5 285.3 209.1 285.9 ;
      RECT  118.7 244.0 119.5 244.8 ;
      RECT  165.5 264.8 166.3 265.6 ;
      RECT  181.3 347.7 181.9 348.3 ;
      RECT  194.9 243.7 195.5 244.3 ;
      RECT  188.0 285.2 188.8 286.0 ;
      RECT  208.5 264.5 209.1 265.1 ;
      RECT  118.7 202.4 119.5 203.2 ;
      RECT  197.2 130.4 198.0 131.2 ;
      RECT  103.7 202.4 104.5 203.2 ;
      RECT  181.3 264.5 181.9 265.1 ;
      RECT  194.9 202.1 195.5 202.7 ;
      RECT  195.6 79.0 196.4 79.8 ;
      RECT  208.5 347.7 209.1 348.3 ;
      RECT  201.7 202.1 202.3 202.7 ;
      RECT  181.3 202.1 181.9 202.7 ;
      RECT  202.4 79.0 203.2 79.8 ;
      RECT  144.7 244.0 145.5 244.8 ;
      RECT  144.7 327.2 145.5 328.0 ;
      RECT  188.0 306.0 188.8 306.8 ;
      RECT  118.7 223.2 119.5 224.0 ;
      RECT  201.7 222.9 202.3 223.5 ;
      RECT  201.7 264.5 202.3 265.1 ;
      RECT  181.3 181.3 181.9 181.9 ;
      RECT  208.5 368.5 209.1 369.1 ;
      RECT  208.5 326.9 209.1 327.5 ;
      RECT  201.4 160.8 202.2 161.6 ;
      RECT  144.7 285.6 145.5 286.4 ;
      RECT  201.7 326.9 202.3 327.5 ;
      RECT  208.5 202.1 209.1 202.7 ;
      RECT  204.0 130.4 204.8 131.2 ;
      RECT  165.5 327.2 166.3 328.0 ;
      RECT  144.7 264.8 145.5 265.6 ;
      RECT  181.3 243.7 181.9 244.3 ;
      RECT  188.0 368.4 188.8 369.2 ;
      RECT  165.5 348.0 166.3 348.8 ;
      RECT  194.6 160.8 195.4 161.6 ;
      RECT  198.2 143.8 199.0 144.6 ;
      RECT  184.6 217.8 185.4 218.6 ;
      RECT  191.5 280.3 192.1 280.9 ;
      RECT  103.7 275.2 104.5 276.0 ;
      RECT  191.4 280.2 192.2 281.0 ;
      RECT  177.9 311.1 178.5 311.7 ;
      RECT  205.1 290.3 205.7 290.9 ;
      RECT  205.0 143.8 205.8 144.6 ;
      RECT  198.3 238.7 198.9 239.3 ;
      RECT  211.9 321.9 212.5 322.5 ;
      RECT  191.4 352.6 192.2 353.4 ;
      RECT  177.9 259.5 178.5 260.1 ;
      RECT  205.1 280.3 205.7 280.9 ;
      RECT  191.4 342.6 192.2 343.4 ;
      RECT  191.5 363.5 192.1 364.1 ;
      RECT  211.9 352.7 212.5 353.3 ;
      RECT  198.3 207.1 198.9 207.7 ;
      RECT  184.7 331.9 185.3 332.5 ;
      RECT  191.4 301.0 192.2 301.8 ;
      RECT  184.7 311.1 185.3 311.7 ;
      RECT  198.3 311.1 198.9 311.7 ;
      RECT  184.7 186.3 185.3 186.9 ;
      RECT  184.7 176.3 185.3 176.9 ;
      RECT  211.9 301.1 212.5 301.7 ;
      RECT  118.7 254.4 119.5 255.2 ;
      RECT  198.3 363.5 198.9 364.1 ;
      RECT  184.7 207.1 185.3 207.7 ;
      RECT  191.4 290.2 192.2 291.0 ;
      RECT  205.1 352.7 205.7 353.3 ;
      RECT  103.7 212.8 104.5 213.6 ;
      RECT  198.3 259.5 198.9 260.1 ;
      RECT  191.5 269.5 192.1 270.1 ;
      RECT  191.5 197.1 192.1 197.7 ;
      RECT  211.9 238.7 212.5 239.3 ;
      RECT  165.5 296.0 166.3 296.8 ;
      RECT  184.7 363.5 185.3 364.1 ;
      RECT  177.9 301.1 178.5 301.7 ;
      RECT  198.3 217.9 198.9 218.5 ;
      RECT  165.5 212.8 166.3 213.6 ;
      RECT  205.1 197.1 205.7 197.7 ;
      RECT  177.9 176.3 178.5 176.9 ;
      RECT  211.9 290.3 212.5 290.9 ;
      RECT  177.9 238.7 178.5 239.3 ;
      RECT  184.6 176.2 185.4 177.0 ;
      RECT  198.3 227.9 198.9 228.5 ;
      RECT  184.7 290.3 185.3 290.9 ;
      RECT  194.2 104.6 195.0 105.4 ;
      RECT  191.5 248.7 192.1 249.3 ;
      RECT  211.9 197.1 212.5 197.7 ;
      RECT  103.7 233.6 104.5 234.4 ;
      RECT  165.5 254.4 166.3 255.2 ;
      RECT  191.5 301.1 192.1 301.7 ;
      RECT  205.1 238.7 205.7 239.3 ;
      RECT  205.1 248.7 205.7 249.3 ;
      RECT  198.3 301.1 198.9 301.7 ;
      RECT  184.6 342.6 185.4 343.4 ;
      RECT  205.1 259.5 205.7 260.1 ;
      RECT  191.5 176.3 192.1 176.9 ;
      RECT  211.9 363.5 212.5 364.1 ;
      RECT  202.4 85.6 203.2 86.4 ;
      RECT  205.1 186.3 205.7 186.9 ;
      RECT  184.6 186.2 185.4 187.0 ;
      RECT  211.9 186.3 212.5 186.9 ;
      RECT  191.4 269.4 192.2 270.2 ;
      RECT  198.3 352.7 198.9 353.3 ;
      RECT  205.1 301.1 205.7 301.7 ;
      RECT  191.5 321.9 192.1 322.5 ;
      RECT  184.7 342.7 185.3 343.3 ;
      RECT  184.6 207.0 185.4 207.8 ;
      RECT  165.5 233.6 166.3 234.4 ;
      RECT  184.7 352.7 185.3 353.3 ;
      RECT  191.5 227.9 192.1 228.5 ;
      RECT  205.1 311.1 205.7 311.7 ;
      RECT  184.6 227.8 185.4 228.6 ;
      RECT  211.9 217.9 212.5 218.5 ;
      RECT  191.5 217.9 192.1 218.5 ;
      RECT  191.4 227.8 192.2 228.6 ;
      RECT  144.7 296.0 145.5 296.8 ;
      RECT  198.3 197.1 198.9 197.7 ;
      RECT  191.4 197.0 192.2 197.8 ;
      RECT  184.7 321.9 185.3 322.5 ;
      RECT  177.9 248.7 178.5 249.3 ;
      RECT  177.9 352.7 178.5 353.3 ;
      RECT  205.1 269.5 205.7 270.1 ;
      RECT  177.9 342.7 178.5 343.3 ;
      RECT  191.5 331.9 192.1 332.5 ;
      RECT  198.3 331.9 198.9 332.5 ;
      RECT  191.4 321.8 192.2 322.6 ;
      RECT  184.6 238.6 185.4 239.4 ;
      RECT  184.6 290.2 185.4 291.0 ;
      RECT  184.7 280.3 185.3 280.9 ;
      RECT  205.1 331.9 205.7 332.5 ;
      RECT  191.4 176.2 192.2 177.0 ;
      RECT  211.9 280.3 212.5 280.9 ;
      RECT  184.7 259.5 185.3 260.1 ;
      RECT  165.5 316.8 166.3 317.6 ;
      RECT  198.3 290.3 198.9 290.9 ;
      RECT  184.6 321.8 185.4 322.6 ;
      RECT  177.9 280.3 178.5 280.9 ;
      RECT  211.9 342.7 212.5 343.3 ;
      RECT  118.7 275.2 119.5 276.0 ;
      RECT  211.9 227.9 212.5 228.5 ;
      RECT  184.6 280.2 185.4 281.0 ;
      RECT  184.7 197.1 185.3 197.7 ;
      RECT  198.3 248.7 198.9 249.3 ;
      RECT  184.7 248.7 185.3 249.3 ;
      RECT  184.6 248.6 185.4 249.4 ;
      RECT  205.1 176.3 205.7 176.9 ;
      RECT  177.9 321.9 178.5 322.5 ;
      RECT  198.3 342.7 198.9 343.3 ;
      RECT  195.6 85.6 196.4 86.4 ;
      RECT  205.1 227.9 205.7 228.5 ;
      RECT  103.7 254.4 104.5 255.2 ;
      RECT  191.4 217.8 192.2 218.6 ;
      RECT  211.9 176.3 212.5 176.9 ;
      RECT  118.7 192.0 119.5 192.8 ;
      RECT  184.6 269.4 185.4 270.2 ;
      RECT  184.7 227.9 185.3 228.5 ;
      RECT  165.5 192.0 166.3 192.8 ;
      RECT  191.5 290.3 192.1 290.9 ;
      RECT  198.3 186.3 198.9 186.9 ;
      RECT  191.5 311.1 192.1 311.7 ;
      RECT  198.3 269.5 198.9 270.1 ;
      RECT  184.6 301.0 185.4 301.8 ;
      RECT  211.9 269.5 212.5 270.1 ;
      RECT  191.4 238.6 192.2 239.4 ;
      RECT  205.1 207.1 205.7 207.7 ;
      RECT  144.7 337.6 145.5 338.4 ;
      RECT  191.5 238.7 192.1 239.3 ;
      RECT  203.8 90.0 204.6 90.8 ;
      RECT  144.7 316.8 145.5 317.6 ;
      RECT  191.4 363.4 192.2 364.2 ;
      RECT  144.7 254.4 145.5 255.2 ;
      RECT  177.9 227.9 178.5 228.5 ;
      RECT  177.9 197.1 178.5 197.7 ;
      RECT  211.9 248.7 212.5 249.3 ;
      RECT  191.4 311.0 192.2 311.8 ;
      RECT  177.9 331.9 178.5 332.5 ;
      RECT  118.7 212.8 119.5 213.6 ;
      RECT  184.7 301.1 185.3 301.7 ;
      RECT  184.6 363.4 185.4 364.2 ;
      RECT  184.6 331.8 185.4 332.6 ;
      RECT  184.6 311.0 185.4 311.8 ;
      RECT  177.9 290.3 178.5 290.9 ;
      RECT  165.5 358.4 166.3 359.2 ;
      RECT  205.1 321.9 205.7 322.5 ;
      RECT  211.9 207.1 212.5 207.7 ;
      RECT  184.7 217.9 185.3 218.5 ;
      RECT  165.5 275.2 166.3 276.0 ;
      RECT  205.1 217.9 205.7 218.5 ;
      RECT  191.4 248.6 192.2 249.4 ;
      RECT  177.9 217.9 178.5 218.5 ;
      RECT  144.7 358.4 145.5 359.2 ;
      RECT  191.5 207.1 192.1 207.7 ;
      RECT  201.0 104.6 201.8 105.4 ;
      RECT  144.7 233.6 145.5 234.4 ;
      RECT  211.9 259.5 212.5 260.1 ;
      RECT  197.0 90.0 197.8 90.8 ;
      RECT  198.3 280.3 198.9 280.9 ;
      RECT  144.7 212.8 145.5 213.6 ;
      RECT  184.6 197.0 185.4 197.8 ;
      RECT  177.9 269.5 178.5 270.1 ;
      RECT  205.1 363.5 205.7 364.1 ;
      RECT  191.5 259.5 192.1 260.1 ;
      RECT  211.9 311.1 212.5 311.7 ;
      RECT  198.3 321.9 198.9 322.5 ;
      RECT  184.7 269.5 185.3 270.1 ;
      RECT  205.1 342.7 205.7 343.3 ;
      RECT  191.4 259.4 192.2 260.2 ;
      RECT  191.4 186.2 192.2 187.0 ;
      RECT  165.5 337.6 166.3 338.4 ;
      RECT  118.7 233.6 119.5 234.4 ;
      RECT  184.7 238.7 185.3 239.3 ;
      RECT  103.7 192.0 104.5 192.8 ;
      RECT  184.6 259.4 185.4 260.2 ;
      RECT  144.7 275.2 145.5 276.0 ;
      RECT  177.9 363.5 178.5 364.1 ;
      RECT  191.5 186.3 192.1 186.9 ;
      RECT  191.5 342.7 192.1 343.3 ;
      RECT  191.5 352.7 192.1 353.3 ;
      RECT  198.3 176.3 198.9 176.9 ;
      RECT  177.9 186.3 178.5 186.9 ;
      RECT  211.9 331.9 212.5 332.5 ;
      RECT  144.7 192.0 145.5 192.8 ;
      RECT  191.4 331.8 192.2 332.6 ;
      RECT  177.9 207.1 178.5 207.7 ;
      RECT  184.6 352.6 185.4 353.4 ;
      RECT  191.4 207.0 192.2 207.8 ;
      RECT  -0.4 19.6 0.4 20.4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
      RECT  -0.4 39.6 0.4 40.4 ;
      RECT  13.2 196.0 12.4 196.8 ;
      RECT  19.6 173.6 18.8 174.4 ;
      RECT  19.6 240.8 18.8 241.6 ;
      RECT  19.6 263.2 18.8 264.0 ;
      RECT  19.6 218.4 18.8 219.2 ;
      RECT  13.2 240.8 12.4 241.6 ;
      RECT  13.2 263.2 12.4 264.0 ;
      RECT  6.8 240.8 6.0 241.6 ;
      RECT  19.6 196.0 18.8 196.8 ;
      RECT  6.8 218.4 6.0 219.2 ;
      RECT  6.8 196.0 6.0 196.8 ;
      RECT  6.8 173.6 6.0 174.4 ;
      RECT  13.2 173.6 12.4 174.4 ;
      RECT  6.8 263.2 6.0 264.0 ;
      RECT  13.2 218.4 12.4 219.2 ;
      RECT  6.8 184.8 6.0 185.6 ;
      RECT  6.8 207.2 6.0 208.0 ;
      RECT  19.6 229.6 18.8 230.4 ;
      RECT  6.8 229.6 6.0 230.4 ;
      RECT  6.8 162.4 6.0 163.2 ;
      RECT  6.8 252.0 6.0 252.8 ;
      RECT  13.2 252.0 12.4 252.8 ;
      RECT  19.6 207.2 18.8 208.0 ;
      RECT  13.2 207.2 12.4 208.0 ;
      RECT  13.2 229.6 12.4 230.4 ;
      RECT  19.6 162.4 18.8 163.2 ;
      RECT  13.2 162.4 12.4 163.2 ;
      RECT  19.6 184.8 18.8 185.6 ;
      RECT  19.6 252.0 18.8 252.8 ;
      RECT  13.2 184.8 12.4 185.6 ;
      RECT  6.0 240.8 6.8 241.6 ;
      RECT  82.6 59.6 83.4 60.4 ;
      RECT  18.8 196.0 19.6 196.8 ;
      RECT  18.8 263.2 19.6 264.0 ;
      RECT  82.6 19.6 83.4 20.4 ;
      RECT  12.4 173.6 13.2 174.4 ;
      RECT  6.0 196.0 6.8 196.8 ;
      RECT  18.8 173.6 19.6 174.4 ;
      RECT  6.0 218.4 6.8 219.2 ;
      RECT  6.0 263.2 6.8 264.0 ;
      RECT  12.4 196.0 13.2 196.8 ;
      RECT  18.8 218.4 19.6 219.2 ;
      RECT  -0.4 19.6 0.4 20.4 ;
      RECT  18.8 240.8 19.6 241.6 ;
      RECT  6.0 173.6 6.8 174.4 ;
      RECT  12.4 263.2 13.2 264.0 ;
      RECT  12.4 218.4 13.2 219.2 ;
      RECT  82.6 139.6 83.4 140.4 ;
      RECT  82.6 99.6 83.4 100.4 ;
      RECT  12.4 240.8 13.2 241.6 ;
      RECT  6.0 229.6 6.8 230.4 ;
      RECT  12.4 207.2 13.2 208.0 ;
      RECT  -0.4 39.6 0.4 40.4 ;
      RECT  12.4 162.4 13.2 163.2 ;
      RECT  82.6 159.6 83.4 160.4 ;
      RECT  82.6 79.6 83.4 80.4 ;
      RECT  12.4 252.0 13.2 252.8 ;
      RECT  82.6 119.6 83.4 120.4 ;
      RECT  18.8 162.4 19.6 163.2 ;
      RECT  12.4 229.6 13.2 230.4 ;
      RECT  18.8 229.6 19.6 230.4 ;
      RECT  82.6 39.6 83.4 40.4 ;
      RECT  6.0 207.2 6.8 208.0 ;
      RECT  6.0 184.8 6.8 185.6 ;
      RECT  18.8 207.2 19.6 208.0 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
      RECT  18.8 252.0 19.6 252.8 ;
      RECT  12.4 184.8 13.2 185.6 ;
      RECT  6.0 252.0 6.8 252.8 ;
      RECT  82.6 -0.4 83.4 0.4 ;
      RECT  18.8 184.8 19.6 185.6 ;
      RECT  6.0 162.4 6.8 163.2 ;
      RECT  62.6 295.7 84.4 296.3 ;
      RECT  73.1 350.2 73.9 351.0 ;
      RECT  73.1 310.2 73.9 311.0 ;
      RECT  73.1 330.2 73.9 331.0 ;
      RECT  73.1 290.2 73.9 291.0 ;
      RECT  73.1 370.2 73.9 371.0 ;
      RECT  178.2 50.9 221.8 51.5 ;
      RECT  188.7 65.4 189.5 66.2 ;
      RECT  210.5 65.4 211.3 66.2 ;
      RECT  188.7 45.4 189.5 46.2 ;
      RECT  210.5 45.4 211.3 46.2 ;
   LAYER  m4 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
